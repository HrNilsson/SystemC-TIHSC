library IEEE;
use IEEE.std_logic_1164.all;  -- defines std_logic types
use IEEE.numeric_std.all;  -- defines add, etc

library UNISIM;
use UNISIM.all; -- defines some Xilinx components, including ROC reset component

use work.craft_gatelibrary.all;
entity SynFir_DoCalculate is 
   port (
      clockin_craft :  in  std_logic;
      syncreset_craft :  in  std_logic;
      asyncreset_craft :  in  std_logic;
      start_craft :  in  std_logic;
      finish_craft :  out  std_logic;
      clock :  in  std_logic;
      reset :  in  std_logic;
      sample_clock :  in  std_logic;
      in_data :  in  std_logic_vector(17 downto 0);
      out_data_out :  out  std_logic_vector(17 downto 0);
      out_data_prev :  in  std_logic_vector(17 downto 0);
      out_data_new :  in  std_logic_vector(17 downto 0);
      in_coef0 :  in  std_logic_vector(31 downto 0);
      in_coef1 :  in  std_logic_vector(31 downto 0);
      in_coef2 :  in  std_logic_vector(31 downto 0);
      in_coef3 :  in  std_logic_vector(31 downto 0);
      in_coef4 :  in  std_logic_vector(31 downto 0);
      in_coef5 :  in  std_logic_vector(31 downto 0);
      in_coef6 :  in  std_logic_vector(31 downto 0);
      in_coef7 :  in  std_logic_vector(31 downto 0);
      in_coef8 :  in  std_logic_vector(31 downto 0);
      in_coef9 :  in  std_logic_vector(31 downto 0);
      in_coef10 :  in  std_logic_vector(31 downto 0);
      in_coef11 :  in  std_logic_vector(31 downto 0);
      in_coef12 :  in  std_logic_vector(31 downto 0);
      in_coef13 :  in  std_logic_vector(31 downto 0);
      in_coef14 :  in  std_logic_vector(31 downto 0);
      in_coef15 :  in  std_logic_vector(31 downto 0);
      in_coef16 :  in  std_logic_vector(31 downto 0);
      in_coef17 :  in  std_logic_vector(31 downto 0);
      in_coef18 :  in  std_logic_vector(31 downto 0);
      in_coef19 :  in  std_logic_vector(31 downto 0);
      in_coef20 :  in  std_logic_vector(31 downto 0);
      in_coef21 :  in  std_logic_vector(31 downto 0);
      in_coef22 :  in  std_logic_vector(31 downto 0);
      m_delay_line_out_0, m_delay_line_out_1, m_delay_line_out_2, m_delay_line_out_3, m_delay_line_out_4, m_delay_line_out_5, m_delay_line_out_6, m_delay_line_out_7, m_delay_line_out_8, m_delay_line_out_9, m_delay_line_out_10, m_delay_line_out_11, m_delay_line_out_12, m_delay_line_out_13, m_delay_line_out_14, m_delay_line_out_15, m_delay_line_out_16, m_delay_line_out_17, m_delay_line_out_18, m_delay_line_out_19, m_delay_line_out_20, m_delay_line_out_21, m_delay_line_out_22 :  out  std_logic_vector(17 downto 0);
      m_delay_line_prev_0, m_delay_line_prev_1, m_delay_line_prev_2, m_delay_line_prev_3, m_delay_line_prev_4, m_delay_line_prev_5, m_delay_line_prev_6, m_delay_line_prev_7, m_delay_line_prev_8, m_delay_line_prev_9, m_delay_line_prev_10, m_delay_line_prev_11, m_delay_line_prev_12, m_delay_line_prev_13, m_delay_line_prev_14, m_delay_line_prev_15, m_delay_line_prev_16, m_delay_line_prev_17, m_delay_line_prev_18, m_delay_line_prev_19, m_delay_line_prev_20, m_delay_line_prev_21, m_delay_line_prev_22 :  in  std_logic_vector(17 downto 0);
      m_delay_line_new_0, m_delay_line_new_1, m_delay_line_new_2, m_delay_line_new_3, m_delay_line_new_4, m_delay_line_new_5, m_delay_line_new_6, m_delay_line_new_7, m_delay_line_new_8, m_delay_line_new_9, m_delay_line_new_10, m_delay_line_new_11, m_delay_line_new_12, m_delay_line_new_13, m_delay_line_new_14, m_delay_line_new_15, m_delay_line_new_16, m_delay_line_new_17, m_delay_line_new_18, m_delay_line_new_19, m_delay_line_new_20, m_delay_line_new_21, m_delay_line_new_22 :  in  std_logic_vector(17 downto 0);
      m_coeffs_out_0, m_coeffs_out_1, m_coeffs_out_2, m_coeffs_out_3, m_coeffs_out_4, m_coeffs_out_5, m_coeffs_out_6, m_coeffs_out_7, m_coeffs_out_8, m_coeffs_out_9, m_coeffs_out_10, m_coeffs_out_11, m_coeffs_out_12, m_coeffs_out_13, m_coeffs_out_14, m_coeffs_out_15, m_coeffs_out_16, m_coeffs_out_17, m_coeffs_out_18, m_coeffs_out_19, m_coeffs_out_20, m_coeffs_out_21, m_coeffs_out_22 :  out  std_logic_vector(31 downto 0);
      m_coeffs_prev_0, m_coeffs_prev_1, m_coeffs_prev_2, m_coeffs_prev_3, m_coeffs_prev_4, m_coeffs_prev_5, m_coeffs_prev_6, m_coeffs_prev_7, m_coeffs_prev_8, m_coeffs_prev_9, m_coeffs_prev_10, m_coeffs_prev_11, m_coeffs_prev_12, m_coeffs_prev_13, m_coeffs_prev_14, m_coeffs_prev_15, m_coeffs_prev_16, m_coeffs_prev_17, m_coeffs_prev_18, m_coeffs_prev_19, m_coeffs_prev_20, m_coeffs_prev_21, m_coeffs_prev_22 :  in  std_logic_vector(31 downto 0);
      m_coeffs_new_0, m_coeffs_new_1, m_coeffs_new_2, m_coeffs_new_3, m_coeffs_new_4, m_coeffs_new_5, m_coeffs_new_6, m_coeffs_new_7, m_coeffs_new_8, m_coeffs_new_9, m_coeffs_new_10, m_coeffs_new_11, m_coeffs_new_12, m_coeffs_new_13, m_coeffs_new_14, m_coeffs_new_15, m_coeffs_new_16, m_coeffs_new_17, m_coeffs_new_18, m_coeffs_new_19, m_coeffs_new_20, m_coeffs_new_21, m_coeffs_new_22 :  in  std_logic_vector(31 downto 0)
   );
end SynFir_DoCalculate;

architecture SynFir_DoCalculate_syn of SynFir_DoCalculate is

   --signal declarations
   signal s0 : std_logic_vector(17 downto 0);
   signal s1_0, s1_1, s1_2, s1_3, s1_4, s1_5, s1_6, s1_7, s1_8, s1_9, s1_10, s1_11, s1_12, s1_13, s1_14, s1_15, s1_16, s1_17, s1_18, s1_19, s1_20, s1_21, s1_22 : std_logic_vector(17 downto 0);
   signal s2_0, s2_1, s2_2, s2_3, s2_4, s2_5, s2_6, s2_7, s2_8, s2_9, s2_10, s2_11, s2_12, s2_13, s2_14, s2_15, s2_16, s2_17, s2_18, s2_19, s2_20, s2_21, s2_22 : std_logic_vector(31 downto 0);
   signal s3 : std_logic;
   signal s4 : std_logic;
   signal s5 : std_logic;
   signal s6 : std_logic;
   signal s7 : std_logic;
   signal s8 : std_logic;
   signal s9 : std_logic;
   signal s10 : std_logic;
   signal s11 : std_logic;
   signal s12 : std_logic;
   signal s13 : std_logic;
   signal s14 : std_logic;
   signal s15 : std_logic_vector(31 downto 0);
   signal s16 : std_logic_vector(31 downto 0);
   signal s17 : std_logic_vector(31 downto 0);
   signal s41 : std_logic;
   signal s19 : std_logic_vector(31 downto 0);
   signal s20 : std_logic_vector(31 downto 0);
   signal s21 : std_logic_vector(31 downto 0);
   signal s22 : std_logic;
   signal s23 : std_logic_vector(31 downto 0);
   signal s24 : std_logic;
   signal s25 : std_logic;
   signal s26 : std_logic_vector(17 downto 0);
   signal s27 : std_logic_vector(4 downto 0);
   signal s28 : std_logic_vector(17 downto 0);
   signal s29 : std_logic_vector(17 downto 0);
   signal s30_0, s30_1, s30_2, s30_3, s30_4, s30_5, s30_6, s30_7, s30_8, s30_9, s30_10, s30_11, s30_12, s30_13, s30_14, s30_15, s30_16, s30_17, s30_18, s30_19, s30_20, s30_21, s30_22 : std_logic_vector(17 downto 0);
   signal s31 : std_logic_vector(31 downto 0);
   signal s32 : std_logic_vector(4 downto 0);
   signal s33 : std_logic_vector(31 downto 0);
   signal s34 : std_logic_vector(31 downto 0);
   signal s35_0, s35_1, s35_2, s35_3, s35_4, s35_5, s35_6, s35_7, s35_8, s35_9, s35_10, s35_11, s35_12, s35_13, s35_14, s35_15, s35_16, s35_17, s35_18, s35_19, s35_20, s35_21, s35_22 : std_logic_vector(31 downto 0);
   signal s36 : std_logic;
   signal s39 : std_logic;
   signal s40 : std_logic;
   signal s42 : std_logic;
   signal s43 : std_logic;
   signal s44 : std_logic;
   signal s45 : std_logic;
   signal s46 : std_logic;
   signal s47 : std_logic;
   signal s48 : std_logic;
   signal s49 : std_logic;
   signal s50 : std_logic;
   signal s51 : std_logic;
   signal s52 : std_logic;
   signal s53 : std_logic;
   signal s54 : std_logic;
   signal s55 : std_logic_vector(31 downto 0);
   signal s56 : std_logic_vector(31 downto 0);
   signal s57 : std_logic_vector(31 downto 0);
   signal s84 : std_logic_vector(17 downto 0);
   signal s59 : std_logic_vector(32 downto 0);
   signal s60 : std_logic_vector(32 downto 0);
   signal s61 : std_logic_vector(32 downto 0);
   signal s62 : std_logic_vector(31 downto 0);
   signal s63 : std_logic_vector(31 downto 0);
   signal s64 : std_logic;
   signal s65 : std_logic_vector(31 downto 0);
   signal s66 : std_logic;
   signal s67 : std_logic;
   signal s68 : std_logic_vector(32 downto 0);
   signal s69 : std_logic_vector(32 downto 0);
   signal s70 : std_logic_vector(32 downto 0);
   signal s71 : std_logic_vector(4 downto 0);
   signal s72 : std_logic_vector(4 downto 0);
   signal s73 : std_logic_vector(17 downto 0);
   signal s74 : std_logic_vector(4 downto 0);
   signal s75 : std_logic_vector(4 downto 0);
   signal s76 : std_logic_vector(17 downto 0);
   signal s77 : std_logic_vector(17 downto 0);
   signal s78_0, s78_1, s78_2, s78_3, s78_4, s78_5, s78_6, s78_7, s78_8, s78_9, s78_10, s78_11, s78_12, s78_13, s78_14, s78_15, s78_16, s78_17, s78_18, s78_19, s78_20, s78_21, s78_22 : std_logic_vector(17 downto 0);
   signal s79 : std_logic;
   signal s82 : std_logic;
   signal s83 : std_logic;
   signal s85 : std_logic_vector(4 downto 0);
   signal s86 : std_logic_vector(17 downto 0);
   signal s87 : std_logic_vector(17 downto 0);
   signal s88_0, s88_1, s88_2, s88_3, s88_4, s88_5, s88_6, s88_7, s88_8, s88_9, s88_10, s88_11, s88_12, s88_13, s88_14, s88_15, s88_16, s88_17, s88_18, s88_19, s88_20, s88_21, s88_22 : std_logic_vector(17 downto 0);
   signal s89 : std_logic_vector(35 downto 0);
   signal s90 : std_logic_vector(35 downto 0);
   signal s91 : std_logic_vector(35 downto 0);
   signal s92 : std_logic_vector(31 downto 0);
   signal s93 : std_logic_vector(31 downto 0);
   signal s94 : std_logic_vector(31 downto 0);
   signal s96 : std_logic_vector(31 downto 0);
   signal s97 : std_logic_vector(31 downto 0);
   signal s98 : std_logic_vector(31 downto 0);
   signal s99 : std_logic;
   signal s100 : std_logic_vector(31 downto 0);
   signal s101 : std_logic;
   signal s102 : std_logic;
   signal s103 : std_logic_vector(64 downto 0);
   signal s104 : std_logic_vector(4 downto 0);
   signal s105 : std_logic_vector(4 downto 0);
   signal s106 : std_logic_vector(17 downto 0);
   signal s107 : std_logic_vector(63 downto 0);
   signal s108 : std_logic_vector(4 downto 0);
   signal s109 : std_logic_vector(4 downto 0);
   signal s110 : std_logic_vector(31 downto 0);
   signal s111 : std_logic_vector(63 downto 0);
   signal s112 : std_logic_vector(63 downto 0);
   signal s113 : std_logic_vector(64 downto 0);
   signal s114 : std_logic_vector(64 downto 0);
   signal s115 : std_logic_vector(35 downto 0);
   signal s116 : std_logic_vector(35 downto 0);
   signal s117 : std_logic;
   signal s120 : std_logic;
   signal s121 : std_logic;
   signal s122 : std_logic_vector(4 downto 0);
   signal s123 : std_logic_vector(35 downto 0);
   signal s124 : std_logic_vector(35 downto 0);
   signal s125 : std_logic_vector(17 downto 0);
   signal s126 : std_logic_vector(17 downto 0);
   signal s127 : std_logic;
   signal s128 : std_logic;
   signal s129 : std_logic;
   signal s130 : std_logic;
   signal s131 : std_logic;
   signal s132 : std_logic;
   signal s133 : std_logic;
   signal s134 : std_logic_vector(31 downto 0);
   signal s135 : std_logic_vector(4 downto 0);
   signal s136 : std_logic_vector(31 downto 0);
   signal s137 : std_logic_vector(31 downto 0);
   signal s138_0, s138_1, s138_2, s138_3, s138_4, s138_5, s138_6, s138_7, s138_8, s138_9, s138_10, s138_11, s138_12, s138_13, s138_14, s138_15, s138_16, s138_17, s138_18, s138_19, s138_20, s138_21, s138_22 : std_logic_vector(31 downto 0);
   signal s139 : std_logic_vector(31 downto 0);
   signal s140 : std_logic_vector(4 downto 0);
   signal s141 : std_logic_vector(31 downto 0);
   signal s142 : std_logic_vector(31 downto 0);
   signal s143_0, s143_1, s143_2, s143_3, s143_4, s143_5, s143_6, s143_7, s143_8, s143_9, s143_10, s143_11, s143_12, s143_13, s143_14, s143_15, s143_16, s143_17, s143_18, s143_19, s143_20, s143_21, s143_22 : std_logic_vector(31 downto 0);
   signal s144 : std_logic_vector(31 downto 0);
   signal s145 : std_logic_vector(4 downto 0);
   signal s146 : std_logic_vector(31 downto 0);
   signal s147 : std_logic_vector(31 downto 0);
   signal s148_0, s148_1, s148_2, s148_3, s148_4, s148_5, s148_6, s148_7, s148_8, s148_9, s148_10, s148_11, s148_12, s148_13, s148_14, s148_15, s148_16, s148_17, s148_18, s148_19, s148_20, s148_21, s148_22 : std_logic_vector(31 downto 0);
   signal s149 : std_logic_vector(31 downto 0);
   signal s150 : std_logic_vector(4 downto 0);
   signal s151 : std_logic_vector(31 downto 0);
   signal s152 : std_logic_vector(31 downto 0);
   signal s153_0, s153_1, s153_2, s153_3, s153_4, s153_5, s153_6, s153_7, s153_8, s153_9, s153_10, s153_11, s153_12, s153_13, s153_14, s153_15, s153_16, s153_17, s153_18, s153_19, s153_20, s153_21, s153_22 : std_logic_vector(31 downto 0);
   signal s154 : std_logic_vector(31 downto 0);
   signal s155 : std_logic_vector(4 downto 0);
   signal s156 : std_logic_vector(31 downto 0);
   signal s157 : std_logic_vector(31 downto 0);
   signal s158_0, s158_1, s158_2, s158_3, s158_4, s158_5, s158_6, s158_7, s158_8, s158_9, s158_10, s158_11, s158_12, s158_13, s158_14, s158_15, s158_16, s158_17, s158_18, s158_19, s158_20, s158_21, s158_22 : std_logic_vector(31 downto 0);
   signal s159 : std_logic_vector(31 downto 0);
   signal s160 : std_logic_vector(4 downto 0);
   signal s161 : std_logic_vector(31 downto 0);
   signal s162 : std_logic_vector(31 downto 0);
   signal s163_0, s163_1, s163_2, s163_3, s163_4, s163_5, s163_6, s163_7, s163_8, s163_9, s163_10, s163_11, s163_12, s163_13, s163_14, s163_15, s163_16, s163_17, s163_18, s163_19, s163_20, s163_21, s163_22 : std_logic_vector(31 downto 0);
   signal s164 : std_logic_vector(31 downto 0);
   signal s165 : std_logic_vector(4 downto 0);
   signal s166 : std_logic_vector(31 downto 0);
   signal s167 : std_logic_vector(31 downto 0);
   signal s168_0, s168_1, s168_2, s168_3, s168_4, s168_5, s168_6, s168_7, s168_8, s168_9, s168_10, s168_11, s168_12, s168_13, s168_14, s168_15, s168_16, s168_17, s168_18, s168_19, s168_20, s168_21, s168_22 : std_logic_vector(31 downto 0);
   signal s169 : std_logic_vector(31 downto 0);
   signal s170 : std_logic_vector(4 downto 0);
   signal s171 : std_logic_vector(31 downto 0);
   signal s172 : std_logic_vector(31 downto 0);
   signal s173_0, s173_1, s173_2, s173_3, s173_4, s173_5, s173_6, s173_7, s173_8, s173_9, s173_10, s173_11, s173_12, s173_13, s173_14, s173_15, s173_16, s173_17, s173_18, s173_19, s173_20, s173_21, s173_22 : std_logic_vector(31 downto 0);
   signal s174 : std_logic_vector(31 downto 0);
   signal s175 : std_logic_vector(4 downto 0);
   signal s176 : std_logic_vector(31 downto 0);
   signal s177 : std_logic_vector(31 downto 0);
   signal s178_0, s178_1, s178_2, s178_3, s178_4, s178_5, s178_6, s178_7, s178_8, s178_9, s178_10, s178_11, s178_12, s178_13, s178_14, s178_15, s178_16, s178_17, s178_18, s178_19, s178_20, s178_21, s178_22 : std_logic_vector(31 downto 0);
   signal s179 : std_logic_vector(31 downto 0);
   signal s180 : std_logic_vector(4 downto 0);
   signal s181 : std_logic_vector(31 downto 0);
   signal s182 : std_logic_vector(31 downto 0);
   signal s183_0, s183_1, s183_2, s183_3, s183_4, s183_5, s183_6, s183_7, s183_8, s183_9, s183_10, s183_11, s183_12, s183_13, s183_14, s183_15, s183_16, s183_17, s183_18, s183_19, s183_20, s183_21, s183_22 : std_logic_vector(31 downto 0);
   signal s184 : std_logic_vector(31 downto 0);
   signal s185 : std_logic_vector(4 downto 0);
   signal s186 : std_logic_vector(31 downto 0);
   signal s187 : std_logic_vector(31 downto 0);
   signal s188_0, s188_1, s188_2, s188_3, s188_4, s188_5, s188_6, s188_7, s188_8, s188_9, s188_10, s188_11, s188_12, s188_13, s188_14, s188_15, s188_16, s188_17, s188_18, s188_19, s188_20, s188_21, s188_22 : std_logic_vector(31 downto 0);
   signal s189 : std_logic_vector(31 downto 0);
   signal s190 : std_logic_vector(4 downto 0);
   signal s191 : std_logic_vector(31 downto 0);
   signal s192 : std_logic_vector(31 downto 0);
   signal s193_0, s193_1, s193_2, s193_3, s193_4, s193_5, s193_6, s193_7, s193_8, s193_9, s193_10, s193_11, s193_12, s193_13, s193_14, s193_15, s193_16, s193_17, s193_18, s193_19, s193_20, s193_21, s193_22 : std_logic_vector(31 downto 0);
   signal s194 : std_logic_vector(31 downto 0);
   signal s195 : std_logic_vector(4 downto 0);
   signal s196 : std_logic_vector(31 downto 0);
   signal s197 : std_logic_vector(31 downto 0);
   signal s198_0, s198_1, s198_2, s198_3, s198_4, s198_5, s198_6, s198_7, s198_8, s198_9, s198_10, s198_11, s198_12, s198_13, s198_14, s198_15, s198_16, s198_17, s198_18, s198_19, s198_20, s198_21, s198_22 : std_logic_vector(31 downto 0);
   signal s199 : std_logic_vector(31 downto 0);
   signal s200 : std_logic_vector(4 downto 0);
   signal s201 : std_logic_vector(31 downto 0);
   signal s202 : std_logic_vector(31 downto 0);
   signal s203_0, s203_1, s203_2, s203_3, s203_4, s203_5, s203_6, s203_7, s203_8, s203_9, s203_10, s203_11, s203_12, s203_13, s203_14, s203_15, s203_16, s203_17, s203_18, s203_19, s203_20, s203_21, s203_22 : std_logic_vector(31 downto 0);
   signal s204 : std_logic_vector(31 downto 0);
   signal s205 : std_logic_vector(4 downto 0);
   signal s206 : std_logic_vector(31 downto 0);
   signal s207 : std_logic_vector(31 downto 0);
   signal s208_0, s208_1, s208_2, s208_3, s208_4, s208_5, s208_6, s208_7, s208_8, s208_9, s208_10, s208_11, s208_12, s208_13, s208_14, s208_15, s208_16, s208_17, s208_18, s208_19, s208_20, s208_21, s208_22 : std_logic_vector(31 downto 0);
   signal s209 : std_logic_vector(31 downto 0);
   signal s210 : std_logic_vector(4 downto 0);
   signal s211 : std_logic_vector(31 downto 0);
   signal s212 : std_logic_vector(31 downto 0);
   signal s213_0, s213_1, s213_2, s213_3, s213_4, s213_5, s213_6, s213_7, s213_8, s213_9, s213_10, s213_11, s213_12, s213_13, s213_14, s213_15, s213_16, s213_17, s213_18, s213_19, s213_20, s213_21, s213_22 : std_logic_vector(31 downto 0);
   signal s214 : std_logic_vector(31 downto 0);
   signal s215 : std_logic_vector(4 downto 0);
   signal s216 : std_logic_vector(31 downto 0);
   signal s217 : std_logic_vector(31 downto 0);
   signal s218_0, s218_1, s218_2, s218_3, s218_4, s218_5, s218_6, s218_7, s218_8, s218_9, s218_10, s218_11, s218_12, s218_13, s218_14, s218_15, s218_16, s218_17, s218_18, s218_19, s218_20, s218_21, s218_22 : std_logic_vector(31 downto 0);
   signal s219 : std_logic_vector(31 downto 0);
   signal s220 : std_logic_vector(4 downto 0);
   signal s221 : std_logic_vector(31 downto 0);
   signal s222 : std_logic_vector(31 downto 0);
   signal s223_0, s223_1, s223_2, s223_3, s223_4, s223_5, s223_6, s223_7, s223_8, s223_9, s223_10, s223_11, s223_12, s223_13, s223_14, s223_15, s223_16, s223_17, s223_18, s223_19, s223_20, s223_21, s223_22 : std_logic_vector(31 downto 0);
   signal s224 : std_logic_vector(31 downto 0);
   signal s225 : std_logic_vector(4 downto 0);
   signal s226 : std_logic_vector(31 downto 0);
   signal s227 : std_logic_vector(31 downto 0);
   signal s228_0, s228_1, s228_2, s228_3, s228_4, s228_5, s228_6, s228_7, s228_8, s228_9, s228_10, s228_11, s228_12, s228_13, s228_14, s228_15, s228_16, s228_17, s228_18, s228_19, s228_20, s228_21, s228_22 : std_logic_vector(31 downto 0);
   signal s229 : std_logic_vector(31 downto 0);
   signal s230 : std_logic_vector(4 downto 0);
   signal s231 : std_logic_vector(31 downto 0);
   signal s232 : std_logic_vector(31 downto 0);
   signal s233_0, s233_1, s233_2, s233_3, s233_4, s233_5, s233_6, s233_7, s233_8, s233_9, s233_10, s233_11, s233_12, s233_13, s233_14, s233_15, s233_16, s233_17, s233_18, s233_19, s233_20, s233_21, s233_22 : std_logic_vector(31 downto 0);
   signal s234 : std_logic_vector(31 downto 0);
   signal s235 : std_logic_vector(4 downto 0);
   signal s236 : std_logic_vector(31 downto 0);
   signal s237 : std_logic_vector(31 downto 0);
   signal s238_0, s238_1, s238_2, s238_3, s238_4, s238_5, s238_6, s238_7, s238_8, s238_9, s238_10, s238_11, s238_12, s238_13, s238_14, s238_15, s238_16, s238_17, s238_18, s238_19, s238_20, s238_21, s238_22 : std_logic_vector(31 downto 0);
   signal s239 : std_logic_vector(31 downto 0);
   signal s240 : std_logic_vector(4 downto 0);
   signal s241 : std_logic_vector(31 downto 0);
   signal s242 : std_logic_vector(31 downto 0);
   signal s243_0, s243_1, s243_2, s243_3, s243_4, s243_5, s243_6, s243_7, s243_8, s243_9, s243_10, s243_11, s243_12, s243_13, s243_14, s243_15, s243_16, s243_17, s243_18, s243_19, s243_20, s243_21, s243_22 : std_logic_vector(31 downto 0);
   signal s244 : std_logic_vector(31 downto 0);
   signal s245 : std_logic_vector(4 downto 0);
   signal s246 : std_logic_vector(31 downto 0);
   signal s247 : std_logic_vector(31 downto 0);
   signal s248_0, s248_1, s248_2, s248_3, s248_4, s248_5, s248_6, s248_7, s248_8, s248_9, s248_10, s248_11, s248_12, s248_13, s248_14, s248_15, s248_16, s248_17, s248_18, s248_19, s248_20, s248_21, s248_22 : std_logic_vector(31 downto 0);
   signal s249 : std_logic;
   signal s250 : std_logic;
   signal s251 : std_logic;
   signal s252 : std_logic;
   signal s253 : std_logic;
   signal s256 : std_logic;
   signal s257 : std_logic;
   signal s302 : std_logic;
   signal s303 : std_logic;
   signal s304 : std_logic;
   signal s305 : std_logic;
   signal s306 : std_logic_vector(4 downto 0);
   signal s309 : std_logic;
   signal s310 : std_logic;
   signal s311 : std_logic;
   signal s312 : std_logic;
   signal s313 : std_logic_vector(4 downto 0);
   signal s316 : std_logic_vector(28 downto 0);
   signal s317 : std_logic_vector(28 downto 0);
   signal s318 : std_logic_vector(28 downto 0);
   signal s319 : std_logic;
   signal s320 : std_logic_vector(5 downto 0);
   signal s323 : std_logic_vector(45 downto 0);
   signal s324 : std_logic_vector(45 downto 0);
   signal s325 : std_logic_vector(45 downto 0);
   signal s326 : std_logic;
   signal s327 : std_logic_vector(4 downto 0);
   signal s330 : std_logic_vector(31 downto 0);
   signal s331 : std_logic_vector(31 downto 0);
   signal s332 : std_logic_vector(31 downto 0);
   signal s333 : std_logic;
   signal s334 : std_logic_vector(4 downto 0);
   signal s337 : std_logic;
   signal s338 : std_logic;
   signal s339 : std_logic;
   signal s340 : std_logic;
   signal s341 : std_logic_vector(5 downto 0);


   --component declarations
   component ROC -- the Xilinx reset component
     port (O : out std_logic);
   end component; --ROC


begin -- body of SynFir_DoCalculate_syn

   -- port connections
   s3 <= clockin_craft;
   s4 <= syncreset_craft;
   s5 <= asyncreset_craft;
   s6 <= start_craft;
   finish_craft <= s257;
   s10 <= reset;
   s46 <= sample_clock;
   s84 <= in_data;
   out_data_out <= s126;
   s0 <= out_data_new;
   s134 <= in_coef0;
   s139 <= in_coef1;
   s144 <= in_coef2;
   s149 <= in_coef3;
   s154 <= in_coef4;
   s159 <= in_coef5;
   s164 <= in_coef6;
   s169 <= in_coef7;
   s174 <= in_coef8;
   s179 <= in_coef9;
   s184 <= in_coef10;
   s189 <= in_coef11;
   s194 <= in_coef12;
   s199 <= in_coef13;
   s204 <= in_coef14;
   s209 <= in_coef15;
   s214 <= in_coef16;
   s219 <= in_coef17;
   s224 <= in_coef18;
   s229 <= in_coef19;
   s234 <= in_coef20;
   s239 <= in_coef21;
   s244 <= in_coef22;
   m_delay_line_out_0 <= s88_0;
   m_delay_line_out_1 <= s88_1;
   m_delay_line_out_2 <= s88_2;
   m_delay_line_out_3 <= s88_3;
   m_delay_line_out_4 <= s88_4;
   m_delay_line_out_5 <= s88_5;
   m_delay_line_out_6 <= s88_6;
   m_delay_line_out_7 <= s88_7;
   m_delay_line_out_8 <= s88_8;
   m_delay_line_out_9 <= s88_9;
   m_delay_line_out_10 <= s88_10;
   m_delay_line_out_11 <= s88_11;
   m_delay_line_out_12 <= s88_12;
   m_delay_line_out_13 <= s88_13;
   m_delay_line_out_14 <= s88_14;
   m_delay_line_out_15 <= s88_15;
   m_delay_line_out_16 <= s88_16;
   m_delay_line_out_17 <= s88_17;
   m_delay_line_out_18 <= s88_18;
   m_delay_line_out_19 <= s88_19;
   m_delay_line_out_20 <= s88_20;
   m_delay_line_out_21 <= s88_21;
   m_delay_line_out_22 <= s88_22;
   s1_0 <= m_delay_line_new_0;
   s1_1 <= m_delay_line_new_1;
   s1_2 <= m_delay_line_new_2;
   s1_3 <= m_delay_line_new_3;
   s1_4 <= m_delay_line_new_4;
   s1_5 <= m_delay_line_new_5;
   s1_6 <= m_delay_line_new_6;
   s1_7 <= m_delay_line_new_7;
   s1_8 <= m_delay_line_new_8;
   s1_9 <= m_delay_line_new_9;
   s1_10 <= m_delay_line_new_10;
   s1_11 <= m_delay_line_new_11;
   s1_12 <= m_delay_line_new_12;
   s1_13 <= m_delay_line_new_13;
   s1_14 <= m_delay_line_new_14;
   s1_15 <= m_delay_line_new_15;
   s1_16 <= m_delay_line_new_16;
   s1_17 <= m_delay_line_new_17;
   s1_18 <= m_delay_line_new_18;
   s1_19 <= m_delay_line_new_19;
   s1_20 <= m_delay_line_new_20;
   s1_21 <= m_delay_line_new_21;
   s1_22 <= m_delay_line_new_22;
   m_coeffs_out_0 <= s248_0;
   m_coeffs_out_1 <= s248_1;
   m_coeffs_out_2 <= s248_2;
   m_coeffs_out_3 <= s248_3;
   m_coeffs_out_4 <= s248_4;
   m_coeffs_out_5 <= s248_5;
   m_coeffs_out_6 <= s248_6;
   m_coeffs_out_7 <= s248_7;
   m_coeffs_out_8 <= s248_8;
   m_coeffs_out_9 <= s248_9;
   m_coeffs_out_10 <= s248_10;
   m_coeffs_out_11 <= s248_11;
   m_coeffs_out_12 <= s248_12;
   m_coeffs_out_13 <= s248_13;
   m_coeffs_out_14 <= s248_14;
   m_coeffs_out_15 <= s248_15;
   m_coeffs_out_16 <= s248_16;
   m_coeffs_out_17 <= s248_17;
   m_coeffs_out_18 <= s248_18;
   m_coeffs_out_19 <= s248_19;
   m_coeffs_out_20 <= s248_20;
   m_coeffs_out_21 <= s248_21;
   m_coeffs_out_22 <= s248_22;
   s2_0 <= m_coeffs_new_0;
   s2_1 <= m_coeffs_new_1;
   s2_2 <= m_coeffs_new_2;
   s2_3 <= m_coeffs_new_3;
   s2_4 <= m_coeffs_new_4;
   s2_5 <= m_coeffs_new_5;
   s2_6 <= m_coeffs_new_6;
   s2_7 <= m_coeffs_new_7;
   s2_8 <= m_coeffs_new_8;
   s2_9 <= m_coeffs_new_9;
   s2_10 <= m_coeffs_new_10;
   s2_11 <= m_coeffs_new_11;
   s2_12 <= m_coeffs_new_12;
   s2_13 <= m_coeffs_new_13;
   s2_14 <= m_coeffs_new_14;
   s2_15 <= m_coeffs_new_15;
   s2_16 <= m_coeffs_new_16;
   s2_17 <= m_coeffs_new_17;
   s2_18 <= m_coeffs_new_18;
   s2_19 <= m_coeffs_new_19;
   s2_20 <= m_coeffs_new_20;
   s2_21 <= m_coeffs_new_21;
   s2_22 <= m_coeffs_new_22;


   s8 <= '1';  -- constint module constint_1_0

   s11 <= s10;  -- ranger typeconverter_1

   s12 <= '1';  -- constint module constint_1_2

   s13 <= equal(s11,s12);  -- relop equal equal_module_3

   s14 <= s13 and s9;  -- and2 and2_4

   s15 <= "00000000000000000000000000000000";  -- constint module constint_0_5

   -- register reg_i_6
   process (s3)
   begin
   if s3'event and s3='1' then  
     s16 <= s21;
   end if;
   end process;

   -- mux2x1 module mux2x1_7
   process(s14, s16, s15)
   begin
   if ( s14 = '1') then s17 <= s15; else s17 <= s16;
   end if;
   end process;

   s19 <= "00000000000000000000000000000001";  -- constint module constint_1_8

   s20 <= to_unsigned(s19) + to_unsigned(s17);  -- add module add_9

   -- mux2x1 module mux2x1_10
   process(s36, s17, s20)
   begin
   if ( s36 = '1') then s21 <= s20; else s21 <= s17;
   end if;
   end process;

   s23 <= "00000000000000000000000000010111";  -- constint module constint_23_11

   s24 <= less_unsigned(s21,s23);  -- relop unsigned less unsigned_less_12

   s26 <= "000000000000000000";  -- constint module constint_0_13

   s27 <= s21(4 downto 0);  -- ranger truncator_14

   -- array reader array_reader_15
   process(s1_0, s1_1, s1_2, s1_3, s1_4, s1_5, s1_6, s1_7, s1_8, s1_9, s1_10, s1_11, s1_12, s1_13, s1_14, s1_15, s1_16, s1_17, s1_18, s1_19, s1_20, s1_21, s1_22, s27)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s27, const00000) = '1' ) then s28 <= s1_0; else
       if (equal(s27, const00001) = '1' ) then s28 <= s1_1; else
       if (equal(s27, const00010) = '1' ) then s28 <= s1_2; else
       if (equal(s27, const00011) = '1' ) then s28 <= s1_3; else
       if (equal(s27, const00100) = '1' ) then s28 <= s1_4; else
       if (equal(s27, const00101) = '1' ) then s28 <= s1_5; else
       if (equal(s27, const00110) = '1' ) then s28 <= s1_6; else
       if (equal(s27, const00111) = '1' ) then s28 <= s1_7; else
       if (equal(s27, const01000) = '1' ) then s28 <= s1_8; else
       if (equal(s27, const01001) = '1' ) then s28 <= s1_9; else
       if (equal(s27, const01010) = '1' ) then s28 <= s1_10; else
       if (equal(s27, const01011) = '1' ) then s28 <= s1_11; else
       if (equal(s27, const01100) = '1' ) then s28 <= s1_12; else
       if (equal(s27, const01101) = '1' ) then s28 <= s1_13; else
       if (equal(s27, const01110) = '1' ) then s28 <= s1_14; else
       if (equal(s27, const01111) = '1' ) then s28 <= s1_15; else
       if (equal(s27, const10000) = '1' ) then s28 <= s1_16; else
       if (equal(s27, const10001) = '1' ) then s28 <= s1_17; else
       if (equal(s27, const10010) = '1' ) then s28 <= s1_18; else
       if (equal(s27, const10011) = '1' ) then s28 <= s1_19; else
       if (equal(s27, const10100) = '1' ) then s28 <= s1_20; else
       if (equal(s27, const10101) = '1' ) then s28 <= s1_21; else
       s28 <= s1_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_16
   process(s25, s28, s26)
   begin
   if ( s25 = '1') then s29 <= s26; else s29 <= s28;
   end if;
   end process;

   -- array writer array_writer_17
   process(s1_0, s1_1, s1_2, s1_3, s1_4, s1_5, s1_6, s1_7, s1_8, s1_9, s1_10, s1_11, s1_12, s1_13, s1_14, s1_15, s1_16, s1_17, s1_18, s1_19, s1_20, s1_21, s1_22, s27, s29)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s27, const00000) = '1' then s30_0 <= s29; else s30_0 <= s1_0; end if;
     if equal(s27, const00001) = '1' then s30_1 <= s29; else s30_1 <= s1_1; end if;
     if equal(s27, const00010) = '1' then s30_2 <= s29; else s30_2 <= s1_2; end if;
     if equal(s27, const00011) = '1' then s30_3 <= s29; else s30_3 <= s1_3; end if;
     if equal(s27, const00100) = '1' then s30_4 <= s29; else s30_4 <= s1_4; end if;
     if equal(s27, const00101) = '1' then s30_5 <= s29; else s30_5 <= s1_5; end if;
     if equal(s27, const00110) = '1' then s30_6 <= s29; else s30_6 <= s1_6; end if;
     if equal(s27, const00111) = '1' then s30_7 <= s29; else s30_7 <= s1_7; end if;
     if equal(s27, const01000) = '1' then s30_8 <= s29; else s30_8 <= s1_8; end if;
     if equal(s27, const01001) = '1' then s30_9 <= s29; else s30_9 <= s1_9; end if;
     if equal(s27, const01010) = '1' then s30_10 <= s29; else s30_10 <= s1_10; end if;
     if equal(s27, const01011) = '1' then s30_11 <= s29; else s30_11 <= s1_11; end if;
     if equal(s27, const01100) = '1' then s30_12 <= s29; else s30_12 <= s1_12; end if;
     if equal(s27, const01101) = '1' then s30_13 <= s29; else s30_13 <= s1_13; end if;
     if equal(s27, const01110) = '1' then s30_14 <= s29; else s30_14 <= s1_14; end if;
     if equal(s27, const01111) = '1' then s30_15 <= s29; else s30_15 <= s1_15; end if;
     if equal(s27, const10000) = '1' then s30_16 <= s29; else s30_16 <= s1_16; end if;
     if equal(s27, const10001) = '1' then s30_17 <= s29; else s30_17 <= s1_17; end if;
     if equal(s27, const10010) = '1' then s30_18 <= s29; else s30_18 <= s1_18; end if;
     if equal(s27, const10011) = '1' then s30_19 <= s29; else s30_19 <= s1_19; end if;
     if equal(s27, const10100) = '1' then s30_20 <= s29; else s30_20 <= s1_20; end if;
     if equal(s27, const10101) = '1' then s30_21 <= s29; else s30_21 <= s1_21; end if;
     if equal(s27, const10110) = '1' then s30_22 <= s29; else s30_22 <= s1_22; end if;
   end process;

   s31 <= "00000000000000000000000000000000";  -- constint module constint_0_18

   s32 <= s21(4 downto 0);  -- ranger truncator_19

   -- array reader array_reader_20
   process(s2_0, s2_1, s2_2, s2_3, s2_4, s2_5, s2_6, s2_7, s2_8, s2_9, s2_10, s2_11, s2_12, s2_13, s2_14, s2_15, s2_16, s2_17, s2_18, s2_19, s2_20, s2_21, s2_22, s32)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s32, const00000) = '1' ) then s33 <= s2_0; else
       if (equal(s32, const00001) = '1' ) then s33 <= s2_1; else
       if (equal(s32, const00010) = '1' ) then s33 <= s2_2; else
       if (equal(s32, const00011) = '1' ) then s33 <= s2_3; else
       if (equal(s32, const00100) = '1' ) then s33 <= s2_4; else
       if (equal(s32, const00101) = '1' ) then s33 <= s2_5; else
       if (equal(s32, const00110) = '1' ) then s33 <= s2_6; else
       if (equal(s32, const00111) = '1' ) then s33 <= s2_7; else
       if (equal(s32, const01000) = '1' ) then s33 <= s2_8; else
       if (equal(s32, const01001) = '1' ) then s33 <= s2_9; else
       if (equal(s32, const01010) = '1' ) then s33 <= s2_10; else
       if (equal(s32, const01011) = '1' ) then s33 <= s2_11; else
       if (equal(s32, const01100) = '1' ) then s33 <= s2_12; else
       if (equal(s32, const01101) = '1' ) then s33 <= s2_13; else
       if (equal(s32, const01110) = '1' ) then s33 <= s2_14; else
       if (equal(s32, const01111) = '1' ) then s33 <= s2_15; else
       if (equal(s32, const10000) = '1' ) then s33 <= s2_16; else
       if (equal(s32, const10001) = '1' ) then s33 <= s2_17; else
       if (equal(s32, const10010) = '1' ) then s33 <= s2_18; else
       if (equal(s32, const10011) = '1' ) then s33 <= s2_19; else
       if (equal(s32, const10100) = '1' ) then s33 <= s2_20; else
       if (equal(s32, const10101) = '1' ) then s33 <= s2_21; else
       s33 <= s2_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_21
   process(s25, s33, s31)
   begin
   if ( s25 = '1') then s34 <= s31; else s34 <= s33;
   end if;
   end process;

   -- array writer array_writer_22
   process(s2_0, s2_1, s2_2, s2_3, s2_4, s2_5, s2_6, s2_7, s2_8, s2_9, s2_10, s2_11, s2_12, s2_13, s2_14, s2_15, s2_16, s2_17, s2_18, s2_19, s2_20, s2_21, s2_22, s32, s34)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s32, const00000) = '1' then s35_0 <= s34; else s35_0 <= s2_0; end if;
     if equal(s32, const00001) = '1' then s35_1 <= s34; else s35_1 <= s2_1; end if;
     if equal(s32, const00010) = '1' then s35_2 <= s34; else s35_2 <= s2_2; end if;
     if equal(s32, const00011) = '1' then s35_3 <= s34; else s35_3 <= s2_3; end if;
     if equal(s32, const00100) = '1' then s35_4 <= s34; else s35_4 <= s2_4; end if;
     if equal(s32, const00101) = '1' then s35_5 <= s34; else s35_5 <= s2_5; end if;
     if equal(s32, const00110) = '1' then s35_6 <= s34; else s35_6 <= s2_6; end if;
     if equal(s32, const00111) = '1' then s35_7 <= s34; else s35_7 <= s2_7; end if;
     if equal(s32, const01000) = '1' then s35_8 <= s34; else s35_8 <= s2_8; end if;
     if equal(s32, const01001) = '1' then s35_9 <= s34; else s35_9 <= s2_9; end if;
     if equal(s32, const01010) = '1' then s35_10 <= s34; else s35_10 <= s2_10; end if;
     if equal(s32, const01011) = '1' then s35_11 <= s34; else s35_11 <= s2_11; end if;
     if equal(s32, const01100) = '1' then s35_12 <= s34; else s35_12 <= s2_12; end if;
     if equal(s32, const01101) = '1' then s35_13 <= s34; else s35_13 <= s2_13; end if;
     if equal(s32, const01110) = '1' then s35_14 <= s34; else s35_14 <= s2_14; end if;
     if equal(s32, const01111) = '1' then s35_15 <= s34; else s35_15 <= s2_15; end if;
     if equal(s32, const10000) = '1' then s35_16 <= s34; else s35_16 <= s2_16; end if;
     if equal(s32, const10001) = '1' then s35_17 <= s34; else s35_17 <= s2_17; end if;
     if equal(s32, const10010) = '1' then s35_18 <= s34; else s35_18 <= s2_18; end if;
     if equal(s32, const10011) = '1' then s35_19 <= s34; else s35_19 <= s2_19; end if;
     if equal(s32, const10100) = '1' then s35_20 <= s34; else s35_20 <= s2_20; end if;
     if equal(s32, const10101) = '1' then s35_21 <= s34; else s35_21 <= s2_21; end if;
     if equal(s32, const10110) = '1' then s35_22 <= s34; else s35_22 <= s2_22; end if;
   end process;

   -- register state_reg_23
   process (s3, s4, s5)
   begin
   if s5 = '1' then
     s36 <= '0';
   elsif s3'event and s3='1' then  
     if s4 = '1' then
        s36 <= '0';
     else
        s36 <= s25;
     end if;
   end if;
   end process;

   s22 <= s14 or s36;  -- or2 or2_24

   s25 <= s22 and s24;  -- and2 and2_25

   s39 <= not s24;  -- not module inv_26

   s40 <= s22 and s39;  -- and2 and2_27

   s41 <= '1';  -- constint module constint_1_28

   -- register reg_clock_state_29
   process (s3)
   begin
   if s3'event and s3='1' then  
     s42 <= s250;
   end if;
   end process;

   -- mux2x1 module mux2x1_30
   process(s40, s42, s41)
   begin
   if ( s40 = '1') then s43 <= s41; else s43 <= s42;
   end if;
   end process;

   s44 <= not s13;  -- not module inv_31

   s45 <= s44 and s9;  -- and2 and2_32

   s47 <= s46;  -- ranger typeconverter_33

   s48 <= '1';  -- constint module constint_1_34

   s49 <= equal(s47,s48);  -- relop equal equal_module_35

   s50 <= s49 and s45;  -- and2 and2_36

   s51 <= s43;  -- ranger typeconverter_37

   s52 <= '0';  -- constint module constint_0_38

   s53 <= equal(s51,s52);  -- relop equal equal_module_39

   s54 <= s53 and s50;  -- and2 and2_40

   s55 <= "00000000000000000000000000010110";  -- constint module constint_22_41

   -- register reg_j_42
   process (s3)
   begin
   if s3'event and s3='1' then  
     s56 <= s63;
   end if;
   end process;

   -- mux2x1 module mux2x1_43
   process(s54, s56, s55)
   begin
   if ( s54 = '1') then s57 <= s55; else s57 <= s56;
   end if;
   end process;

   s60 <= "000000000000000000000000000000001";  -- constint module constint_1_45

   s61 <= to_unsigned(s59) - to_unsigned(s60);  -- minus module sub_46

   s62 <= s61(31 downto 0);  -- ranger truncator_47

   -- mux2x1 module mux2x1_48
   process(s79, s57, s62)
   begin
   if ( s79 = '1') then s63 <= s62; else s63 <= s57;
   end if;
   end process;

   s65 <= "00000000000000000000000000000000";  -- constint module constint_0_49

   s66 <= greater_signed(s63,s65);  -- relop signed greater signed_greater_50

   s69 <= "000000000000000000000000000000001";  -- constint module constint_1_52

   s70 <= to_unsigned(s68) - to_unsigned(s69);  -- minus module sub_53

   s71 <= s70(4 downto 0);  -- ranger truncator_54

   s72 <= s71(4 downto 0);  -- ranger typeconverter_55

   -- array reader array_reader_56
   process(s30_0, s30_1, s30_2, s30_3, s30_4, s30_5, s30_6, s30_7, s30_8, s30_9, s30_10, s30_11, s30_12, s30_13, s30_14, s30_15, s30_16, s30_17, s30_18, s30_19, s30_20, s30_21, s30_22, s72)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s72, const00000) = '1' ) then s73 <= s30_0; else
       if (equal(s72, const00001) = '1' ) then s73 <= s30_1; else
       if (equal(s72, const00010) = '1' ) then s73 <= s30_2; else
       if (equal(s72, const00011) = '1' ) then s73 <= s30_3; else
       if (equal(s72, const00100) = '1' ) then s73 <= s30_4; else
       if (equal(s72, const00101) = '1' ) then s73 <= s30_5; else
       if (equal(s72, const00110) = '1' ) then s73 <= s30_6; else
       if (equal(s72, const00111) = '1' ) then s73 <= s30_7; else
       if (equal(s72, const01000) = '1' ) then s73 <= s30_8; else
       if (equal(s72, const01001) = '1' ) then s73 <= s30_9; else
       if (equal(s72, const01010) = '1' ) then s73 <= s30_10; else
       if (equal(s72, const01011) = '1' ) then s73 <= s30_11; else
       if (equal(s72, const01100) = '1' ) then s73 <= s30_12; else
       if (equal(s72, const01101) = '1' ) then s73 <= s30_13; else
       if (equal(s72, const01110) = '1' ) then s73 <= s30_14; else
       if (equal(s72, const01111) = '1' ) then s73 <= s30_15; else
       if (equal(s72, const10000) = '1' ) then s73 <= s30_16; else
       if (equal(s72, const10001) = '1' ) then s73 <= s30_17; else
       if (equal(s72, const10010) = '1' ) then s73 <= s30_18; else
       if (equal(s72, const10011) = '1' ) then s73 <= s30_19; else
       if (equal(s72, const10100) = '1' ) then s73 <= s30_20; else
       if (equal(s72, const10101) = '1' ) then s73 <= s30_21; else
       s73 <= s30_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   s74 <= s63(4 downto 0);  -- ranger truncator_57

   s75 <= s74(4 downto 0);  -- ranger typeconverter_58

   -- array reader array_reader_59
   process(s30_0, s30_1, s30_2, s30_3, s30_4, s30_5, s30_6, s30_7, s30_8, s30_9, s30_10, s30_11, s30_12, s30_13, s30_14, s30_15, s30_16, s30_17, s30_18, s30_19, s30_20, s30_21, s30_22, s75)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s75, const00000) = '1' ) then s76 <= s30_0; else
       if (equal(s75, const00001) = '1' ) then s76 <= s30_1; else
       if (equal(s75, const00010) = '1' ) then s76 <= s30_2; else
       if (equal(s75, const00011) = '1' ) then s76 <= s30_3; else
       if (equal(s75, const00100) = '1' ) then s76 <= s30_4; else
       if (equal(s75, const00101) = '1' ) then s76 <= s30_5; else
       if (equal(s75, const00110) = '1' ) then s76 <= s30_6; else
       if (equal(s75, const00111) = '1' ) then s76 <= s30_7; else
       if (equal(s75, const01000) = '1' ) then s76 <= s30_8; else
       if (equal(s75, const01001) = '1' ) then s76 <= s30_9; else
       if (equal(s75, const01010) = '1' ) then s76 <= s30_10; else
       if (equal(s75, const01011) = '1' ) then s76 <= s30_11; else
       if (equal(s75, const01100) = '1' ) then s76 <= s30_12; else
       if (equal(s75, const01101) = '1' ) then s76 <= s30_13; else
       if (equal(s75, const01110) = '1' ) then s76 <= s30_14; else
       if (equal(s75, const01111) = '1' ) then s76 <= s30_15; else
       if (equal(s75, const10000) = '1' ) then s76 <= s30_16; else
       if (equal(s75, const10001) = '1' ) then s76 <= s30_17; else
       if (equal(s75, const10010) = '1' ) then s76 <= s30_18; else
       if (equal(s75, const10011) = '1' ) then s76 <= s30_19; else
       if (equal(s75, const10100) = '1' ) then s76 <= s30_20; else
       if (equal(s75, const10101) = '1' ) then s76 <= s30_21; else
       s76 <= s30_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_60
   process(s67, s76, s73)
   begin
   if ( s67 = '1') then s77 <= s73; else s77 <= s76;
   end if;
   end process;

   -- array writer array_writer_61
   process(s30_0, s30_1, s30_2, s30_3, s30_4, s30_5, s30_6, s30_7, s30_8, s30_9, s30_10, s30_11, s30_12, s30_13, s30_14, s30_15, s30_16, s30_17, s30_18, s30_19, s30_20, s30_21, s30_22, s75, s77)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s75, const00000) = '1' then s78_0 <= s77; else s78_0 <= s30_0; end if;
     if equal(s75, const00001) = '1' then s78_1 <= s77; else s78_1 <= s30_1; end if;
     if equal(s75, const00010) = '1' then s78_2 <= s77; else s78_2 <= s30_2; end if;
     if equal(s75, const00011) = '1' then s78_3 <= s77; else s78_3 <= s30_3; end if;
     if equal(s75, const00100) = '1' then s78_4 <= s77; else s78_4 <= s30_4; end if;
     if equal(s75, const00101) = '1' then s78_5 <= s77; else s78_5 <= s30_5; end if;
     if equal(s75, const00110) = '1' then s78_6 <= s77; else s78_6 <= s30_6; end if;
     if equal(s75, const00111) = '1' then s78_7 <= s77; else s78_7 <= s30_7; end if;
     if equal(s75, const01000) = '1' then s78_8 <= s77; else s78_8 <= s30_8; end if;
     if equal(s75, const01001) = '1' then s78_9 <= s77; else s78_9 <= s30_9; end if;
     if equal(s75, const01010) = '1' then s78_10 <= s77; else s78_10 <= s30_10; end if;
     if equal(s75, const01011) = '1' then s78_11 <= s77; else s78_11 <= s30_11; end if;
     if equal(s75, const01100) = '1' then s78_12 <= s77; else s78_12 <= s30_12; end if;
     if equal(s75, const01101) = '1' then s78_13 <= s77; else s78_13 <= s30_13; end if;
     if equal(s75, const01110) = '1' then s78_14 <= s77; else s78_14 <= s30_14; end if;
     if equal(s75, const01111) = '1' then s78_15 <= s77; else s78_15 <= s30_15; end if;
     if equal(s75, const10000) = '1' then s78_16 <= s77; else s78_16 <= s30_16; end if;
     if equal(s75, const10001) = '1' then s78_17 <= s77; else s78_17 <= s30_17; end if;
     if equal(s75, const10010) = '1' then s78_18 <= s77; else s78_18 <= s30_18; end if;
     if equal(s75, const10011) = '1' then s78_19 <= s77; else s78_19 <= s30_19; end if;
     if equal(s75, const10100) = '1' then s78_20 <= s77; else s78_20 <= s30_20; end if;
     if equal(s75, const10101) = '1' then s78_21 <= s77; else s78_21 <= s30_21; end if;
     if equal(s75, const10110) = '1' then s78_22 <= s77; else s78_22 <= s30_22; end if;
   end process;

   -- register state_reg_62
   process (s3, s4, s5)
   begin
   if s5 = '1' then
     s79 <= '0';
   elsif s3'event and s3='1' then  
     if s4 = '1' then
        s79 <= '0';
     else
        s79 <= s67;
     end if;
   end if;
   end process;

   s64 <= s54 or s79;  -- or2 or2_63

   s67 <= s64 and s66;  -- and2 and2_64

   s82 <= not s66;  -- not module inv_65

   s83 <= s64 and s82;  -- and2 and2_66

   s85 <= "00000";  -- constint module constint_0_67

   -- array reader array_reader_68
   process(s78_0, s78_1, s78_2, s78_3, s78_4, s78_5, s78_6, s78_7, s78_8, s78_9, s78_10, s78_11, s78_12, s78_13, s78_14, s78_15, s78_16, s78_17, s78_18, s78_19, s78_20, s78_21, s78_22, s85)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s85, const00000) = '1' ) then s86 <= s78_0; else
       if (equal(s85, const00001) = '1' ) then s86 <= s78_1; else
       if (equal(s85, const00010) = '1' ) then s86 <= s78_2; else
       if (equal(s85, const00011) = '1' ) then s86 <= s78_3; else
       if (equal(s85, const00100) = '1' ) then s86 <= s78_4; else
       if (equal(s85, const00101) = '1' ) then s86 <= s78_5; else
       if (equal(s85, const00110) = '1' ) then s86 <= s78_6; else
       if (equal(s85, const00111) = '1' ) then s86 <= s78_7; else
       if (equal(s85, const01000) = '1' ) then s86 <= s78_8; else
       if (equal(s85, const01001) = '1' ) then s86 <= s78_9; else
       if (equal(s85, const01010) = '1' ) then s86 <= s78_10; else
       if (equal(s85, const01011) = '1' ) then s86 <= s78_11; else
       if (equal(s85, const01100) = '1' ) then s86 <= s78_12; else
       if (equal(s85, const01101) = '1' ) then s86 <= s78_13; else
       if (equal(s85, const01110) = '1' ) then s86 <= s78_14; else
       if (equal(s85, const01111) = '1' ) then s86 <= s78_15; else
       if (equal(s85, const10000) = '1' ) then s86 <= s78_16; else
       if (equal(s85, const10001) = '1' ) then s86 <= s78_17; else
       if (equal(s85, const10010) = '1' ) then s86 <= s78_18; else
       if (equal(s85, const10011) = '1' ) then s86 <= s78_19; else
       if (equal(s85, const10100) = '1' ) then s86 <= s78_20; else
       if (equal(s85, const10101) = '1' ) then s86 <= s78_21; else
       s86 <= s78_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_69
   process(s83, s86, s84)
   begin
   if ( s83 = '1') then s87 <= s84; else s87 <= s86;
   end if;
   end process;

   -- array writer array_writer_70
   process(s78_0, s78_1, s78_2, s78_3, s78_4, s78_5, s78_6, s78_7, s78_8, s78_9, s78_10, s78_11, s78_12, s78_13, s78_14, s78_15, s78_16, s78_17, s78_18, s78_19, s78_20, s78_21, s78_22, s85, s87)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s85, const00000) = '1' then s88_0 <= s87; else s88_0 <= s78_0; end if;
     if equal(s85, const00001) = '1' then s88_1 <= s87; else s88_1 <= s78_1; end if;
     if equal(s85, const00010) = '1' then s88_2 <= s87; else s88_2 <= s78_2; end if;
     if equal(s85, const00011) = '1' then s88_3 <= s87; else s88_3 <= s78_3; end if;
     if equal(s85, const00100) = '1' then s88_4 <= s87; else s88_4 <= s78_4; end if;
     if equal(s85, const00101) = '1' then s88_5 <= s87; else s88_5 <= s78_5; end if;
     if equal(s85, const00110) = '1' then s88_6 <= s87; else s88_6 <= s78_6; end if;
     if equal(s85, const00111) = '1' then s88_7 <= s87; else s88_7 <= s78_7; end if;
     if equal(s85, const01000) = '1' then s88_8 <= s87; else s88_8 <= s78_8; end if;
     if equal(s85, const01001) = '1' then s88_9 <= s87; else s88_9 <= s78_9; end if;
     if equal(s85, const01010) = '1' then s88_10 <= s87; else s88_10 <= s78_10; end if;
     if equal(s85, const01011) = '1' then s88_11 <= s87; else s88_11 <= s78_11; end if;
     if equal(s85, const01100) = '1' then s88_12 <= s87; else s88_12 <= s78_12; end if;
     if equal(s85, const01101) = '1' then s88_13 <= s87; else s88_13 <= s78_13; end if;
     if equal(s85, const01110) = '1' then s88_14 <= s87; else s88_14 <= s78_14; end if;
     if equal(s85, const01111) = '1' then s88_15 <= s87; else s88_15 <= s78_15; end if;
     if equal(s85, const10000) = '1' then s88_16 <= s87; else s88_16 <= s78_16; end if;
     if equal(s85, const10001) = '1' then s88_17 <= s87; else s88_17 <= s78_17; end if;
     if equal(s85, const10010) = '1' then s88_18 <= s87; else s88_18 <= s78_18; end if;
     if equal(s85, const10011) = '1' then s88_19 <= s87; else s88_19 <= s78_19; end if;
     if equal(s85, const10100) = '1' then s88_20 <= s87; else s88_20 <= s78_20; end if;
     if equal(s85, const10101) = '1' then s88_21 <= s87; else s88_21 <= s78_21; end if;
     if equal(s85, const10110) = '1' then s88_22 <= s87; else s88_22 <= s78_22; end if;
   end process;

   s89 <= "000000000000000000000000000000000000";  -- constint module constint_0_71

   -- register reg_sum_72
   process (s3)
   begin
   if s3'event and s3='1' then  
     s90 <= s124;
   end if;
   end process;

   -- mux2x1 module mux2x1_73
   process(s83, s90, s89)
   begin
   if ( s83 = '1') then s91 <= s89; else s91 <= s90;
   end if;
   end process;

   s92 <= "00000000000000000000000000000000";  -- constint module constint_0_74

   -- register reg_i_75
   process (s3)
   begin
   if s3'event and s3='1' then  
     s93 <= s98;
   end if;
   end process;

   -- mux2x1 module mux2x1_76
   process(s83, s93, s92)
   begin
   if ( s83 = '1') then s94 <= s92; else s94 <= s93;
   end if;
   end process;

   s96 <= "00000000000000000000000000000001";  -- constint module constint_1_77

   s97 <= to_unsigned(s96) + to_unsigned(s94);  -- add module add_78

   -- mux2x1 module mux2x1_79
   process(s117, s94, s97)
   begin
   if ( s117 = '1') then s98 <= s97; else s98 <= s94;
   end if;
   end process;

   s100 <= "00000000000000000000000000010111";  -- constint module constint_23_80

   s101 <= less_signed(s98,s100);  -- relop signed less signed_less_81

   s104 <= s98(4 downto 0);  -- ranger truncator_83

   s105 <= s104(4 downto 0);  -- ranger typeconverter_84

   -- array reader array_reader_85
   process(s88_0, s88_1, s88_2, s88_3, s88_4, s88_5, s88_6, s88_7, s88_8, s88_9, s88_10, s88_11, s88_12, s88_13, s88_14, s88_15, s88_16, s88_17, s88_18, s88_19, s88_20, s88_21, s88_22, s105)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s105, const00000) = '1' ) then s106 <= s88_0; else
       if (equal(s105, const00001) = '1' ) then s106 <= s88_1; else
       if (equal(s105, const00010) = '1' ) then s106 <= s88_2; else
       if (equal(s105, const00011) = '1' ) then s106 <= s88_3; else
       if (equal(s105, const00100) = '1' ) then s106 <= s88_4; else
       if (equal(s105, const00101) = '1' ) then s106 <= s88_5; else
       if (equal(s105, const00110) = '1' ) then s106 <= s88_6; else
       if (equal(s105, const00111) = '1' ) then s106 <= s88_7; else
       if (equal(s105, const01000) = '1' ) then s106 <= s88_8; else
       if (equal(s105, const01001) = '1' ) then s106 <= s88_9; else
       if (equal(s105, const01010) = '1' ) then s106 <= s88_10; else
       if (equal(s105, const01011) = '1' ) then s106 <= s88_11; else
       if (equal(s105, const01100) = '1' ) then s106 <= s88_12; else
       if (equal(s105, const01101) = '1' ) then s106 <= s88_13; else
       if (equal(s105, const01110) = '1' ) then s106 <= s88_14; else
       if (equal(s105, const01111) = '1' ) then s106 <= s88_15; else
       if (equal(s105, const10000) = '1' ) then s106 <= s88_16; else
       if (equal(s105, const10001) = '1' ) then s106 <= s88_17; else
       if (equal(s105, const10010) = '1' ) then s106 <= s88_18; else
       if (equal(s105, const10011) = '1' ) then s106 <= s88_19; else
       if (equal(s105, const10100) = '1' ) then s106 <= s88_20; else
       if (equal(s105, const10101) = '1' ) then s106 <= s88_21; else
       s106 <= s88_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   s108 <= s98(4 downto 0);  -- ranger truncator_87

   s109 <= s108(4 downto 0);  -- ranger typeconverter_88

   -- array reader array_reader_89
   process(s35_0, s35_1, s35_2, s35_3, s35_4, s35_5, s35_6, s35_7, s35_8, s35_9, s35_10, s35_11, s35_12, s35_13, s35_14, s35_15, s35_16, s35_17, s35_18, s35_19, s35_20, s35_21, s35_22, s109)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s109, const00000) = '1' ) then s110 <= s35_0; else
       if (equal(s109, const00001) = '1' ) then s110 <= s35_1; else
       if (equal(s109, const00010) = '1' ) then s110 <= s35_2; else
       if (equal(s109, const00011) = '1' ) then s110 <= s35_3; else
       if (equal(s109, const00100) = '1' ) then s110 <= s35_4; else
       if (equal(s109, const00101) = '1' ) then s110 <= s35_5; else
       if (equal(s109, const00110) = '1' ) then s110 <= s35_6; else
       if (equal(s109, const00111) = '1' ) then s110 <= s35_7; else
       if (equal(s109, const01000) = '1' ) then s110 <= s35_8; else
       if (equal(s109, const01001) = '1' ) then s110 <= s35_9; else
       if (equal(s109, const01010) = '1' ) then s110 <= s35_10; else
       if (equal(s109, const01011) = '1' ) then s110 <= s35_11; else
       if (equal(s109, const01100) = '1' ) then s110 <= s35_12; else
       if (equal(s109, const01101) = '1' ) then s110 <= s35_13; else
       if (equal(s109, const01110) = '1' ) then s110 <= s35_14; else
       if (equal(s109, const01111) = '1' ) then s110 <= s35_15; else
       if (equal(s109, const10000) = '1' ) then s110 <= s35_16; else
       if (equal(s109, const10001) = '1' ) then s110 <= s35_17; else
       if (equal(s109, const10010) = '1' ) then s110 <= s35_18; else
       if (equal(s109, const10011) = '1' ) then s110 <= s35_19; else
       if (equal(s109, const10100) = '1' ) then s110 <= s35_20; else
       if (equal(s109, const10101) = '1' ) then s110 <= s35_21; else
       s110 <= s35_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   s112 <= to_signed(s107) * to_signed(s111);  -- times signed_mult_91

   s114 <= to_unsigned(s103) + to_unsigned(s113);  -- add module add_93

   s115 <= s114(35 downto 0);  -- ranger truncator_94

   -- mux2x1 module mux2x1_95
   process(s102, s91, s115)
   begin
   if ( s102 = '1') then s116 <= s115; else s116 <= s91;
   end if;
   end process;

   -- register state_reg_96
   process (s3, s4, s5)
   begin
   if s5 = '1' then
     s117 <= '0';
   elsif s3'event and s3='1' then  
     if s4 = '1' then
        s117 <= '0';
     else
        s117 <= s102;
     end if;
   end if;
   end process;

   s99 <= s83 or s117;  -- or2 or2_97

   s102 <= s99 and s101;  -- and2 and2_98

   s120 <= not s101;  -- not module inv_99

   s121 <= s99 and s120;  -- and2 and2_100

   s122 <= "10001";  -- constint module constint_17_101

   -- arithmetic rightshift module arithrightshift_102
   s123 <= to_stdlogicvector(to_bitvector(s116) sra to_integer(to_unsigned(s122)));

   -- mux2x1 module mux2x1_103
   process(s121, s116, s123)
   begin
   if ( s121 = '1') then s124 <= s123; else s124 <= s116;
   end if;
   end process;

   s125 <= s124(17 downto 0);  -- ranger truncator_104

   -- mux2x1 module mux2x1_105
   process(s121, s0, s125)
   begin
   if ( s121 = '1') then s126 <= s125; else s126 <= s0;
   end if;
   end process;

   s127 <= '1';  -- constint module constint_1_106

   -- mux2x1 module mux2x1_107
   process(s121, s43, s127)
   begin
   if ( s121 = '1') then s128 <= s127; else s128 <= s43;
   end if;
   end process;

   s129 <= not s53;  -- not module inv_108

   s130 <= s50 and s129;  -- and2 and2_109

   s131 <= s130 or s121;  -- or2 or2_110

   s132 <= not s49;  -- not module inv_111

   s133 <= s132 and s45;  -- and2 and2_112

   s135 <= "00000";  -- constint module constint_0_113

   -- array reader array_reader_114
   process(s35_0, s35_1, s35_2, s35_3, s35_4, s35_5, s35_6, s35_7, s35_8, s35_9, s35_10, s35_11, s35_12, s35_13, s35_14, s35_15, s35_16, s35_17, s35_18, s35_19, s35_20, s35_21, s35_22, s135)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s135, const00000) = '1' ) then s136 <= s35_0; else
       if (equal(s135, const00001) = '1' ) then s136 <= s35_1; else
       if (equal(s135, const00010) = '1' ) then s136 <= s35_2; else
       if (equal(s135, const00011) = '1' ) then s136 <= s35_3; else
       if (equal(s135, const00100) = '1' ) then s136 <= s35_4; else
       if (equal(s135, const00101) = '1' ) then s136 <= s35_5; else
       if (equal(s135, const00110) = '1' ) then s136 <= s35_6; else
       if (equal(s135, const00111) = '1' ) then s136 <= s35_7; else
       if (equal(s135, const01000) = '1' ) then s136 <= s35_8; else
       if (equal(s135, const01001) = '1' ) then s136 <= s35_9; else
       if (equal(s135, const01010) = '1' ) then s136 <= s35_10; else
       if (equal(s135, const01011) = '1' ) then s136 <= s35_11; else
       if (equal(s135, const01100) = '1' ) then s136 <= s35_12; else
       if (equal(s135, const01101) = '1' ) then s136 <= s35_13; else
       if (equal(s135, const01110) = '1' ) then s136 <= s35_14; else
       if (equal(s135, const01111) = '1' ) then s136 <= s35_15; else
       if (equal(s135, const10000) = '1' ) then s136 <= s35_16; else
       if (equal(s135, const10001) = '1' ) then s136 <= s35_17; else
       if (equal(s135, const10010) = '1' ) then s136 <= s35_18; else
       if (equal(s135, const10011) = '1' ) then s136 <= s35_19; else
       if (equal(s135, const10100) = '1' ) then s136 <= s35_20; else
       if (equal(s135, const10101) = '1' ) then s136 <= s35_21; else
       s136 <= s35_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_115
   process(s133, s136, s134)
   begin
   if ( s133 = '1') then s137 <= s134; else s137 <= s136;
   end if;
   end process;

   -- array writer array_writer_116
   process(s35_0, s35_1, s35_2, s35_3, s35_4, s35_5, s35_6, s35_7, s35_8, s35_9, s35_10, s35_11, s35_12, s35_13, s35_14, s35_15, s35_16, s35_17, s35_18, s35_19, s35_20, s35_21, s35_22, s135, s137)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s135, const00000) = '1' then s138_0 <= s137; else s138_0 <= s35_0; end if;
     if equal(s135, const00001) = '1' then s138_1 <= s137; else s138_1 <= s35_1; end if;
     if equal(s135, const00010) = '1' then s138_2 <= s137; else s138_2 <= s35_2; end if;
     if equal(s135, const00011) = '1' then s138_3 <= s137; else s138_3 <= s35_3; end if;
     if equal(s135, const00100) = '1' then s138_4 <= s137; else s138_4 <= s35_4; end if;
     if equal(s135, const00101) = '1' then s138_5 <= s137; else s138_5 <= s35_5; end if;
     if equal(s135, const00110) = '1' then s138_6 <= s137; else s138_6 <= s35_6; end if;
     if equal(s135, const00111) = '1' then s138_7 <= s137; else s138_7 <= s35_7; end if;
     if equal(s135, const01000) = '1' then s138_8 <= s137; else s138_8 <= s35_8; end if;
     if equal(s135, const01001) = '1' then s138_9 <= s137; else s138_9 <= s35_9; end if;
     if equal(s135, const01010) = '1' then s138_10 <= s137; else s138_10 <= s35_10; end if;
     if equal(s135, const01011) = '1' then s138_11 <= s137; else s138_11 <= s35_11; end if;
     if equal(s135, const01100) = '1' then s138_12 <= s137; else s138_12 <= s35_12; end if;
     if equal(s135, const01101) = '1' then s138_13 <= s137; else s138_13 <= s35_13; end if;
     if equal(s135, const01110) = '1' then s138_14 <= s137; else s138_14 <= s35_14; end if;
     if equal(s135, const01111) = '1' then s138_15 <= s137; else s138_15 <= s35_15; end if;
     if equal(s135, const10000) = '1' then s138_16 <= s137; else s138_16 <= s35_16; end if;
     if equal(s135, const10001) = '1' then s138_17 <= s137; else s138_17 <= s35_17; end if;
     if equal(s135, const10010) = '1' then s138_18 <= s137; else s138_18 <= s35_18; end if;
     if equal(s135, const10011) = '1' then s138_19 <= s137; else s138_19 <= s35_19; end if;
     if equal(s135, const10100) = '1' then s138_20 <= s137; else s138_20 <= s35_20; end if;
     if equal(s135, const10101) = '1' then s138_21 <= s137; else s138_21 <= s35_21; end if;
     if equal(s135, const10110) = '1' then s138_22 <= s137; else s138_22 <= s35_22; end if;
   end process;

   s140 <= "00001";  -- constint module constint_1_117

   -- array reader array_reader_118
   process(s138_0, s138_1, s138_2, s138_3, s138_4, s138_5, s138_6, s138_7, s138_8, s138_9, s138_10, s138_11, s138_12, s138_13, s138_14, s138_15, s138_16, s138_17, s138_18, s138_19, s138_20, s138_21, s138_22, s140)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s140, const00000) = '1' ) then s141 <= s138_0; else
       if (equal(s140, const00001) = '1' ) then s141 <= s138_1; else
       if (equal(s140, const00010) = '1' ) then s141 <= s138_2; else
       if (equal(s140, const00011) = '1' ) then s141 <= s138_3; else
       if (equal(s140, const00100) = '1' ) then s141 <= s138_4; else
       if (equal(s140, const00101) = '1' ) then s141 <= s138_5; else
       if (equal(s140, const00110) = '1' ) then s141 <= s138_6; else
       if (equal(s140, const00111) = '1' ) then s141 <= s138_7; else
       if (equal(s140, const01000) = '1' ) then s141 <= s138_8; else
       if (equal(s140, const01001) = '1' ) then s141 <= s138_9; else
       if (equal(s140, const01010) = '1' ) then s141 <= s138_10; else
       if (equal(s140, const01011) = '1' ) then s141 <= s138_11; else
       if (equal(s140, const01100) = '1' ) then s141 <= s138_12; else
       if (equal(s140, const01101) = '1' ) then s141 <= s138_13; else
       if (equal(s140, const01110) = '1' ) then s141 <= s138_14; else
       if (equal(s140, const01111) = '1' ) then s141 <= s138_15; else
       if (equal(s140, const10000) = '1' ) then s141 <= s138_16; else
       if (equal(s140, const10001) = '1' ) then s141 <= s138_17; else
       if (equal(s140, const10010) = '1' ) then s141 <= s138_18; else
       if (equal(s140, const10011) = '1' ) then s141 <= s138_19; else
       if (equal(s140, const10100) = '1' ) then s141 <= s138_20; else
       if (equal(s140, const10101) = '1' ) then s141 <= s138_21; else
       s141 <= s138_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_119
   process(s133, s141, s139)
   begin
   if ( s133 = '1') then s142 <= s139; else s142 <= s141;
   end if;
   end process;

   -- array writer array_writer_120
   process(s138_0, s138_1, s138_2, s138_3, s138_4, s138_5, s138_6, s138_7, s138_8, s138_9, s138_10, s138_11, s138_12, s138_13, s138_14, s138_15, s138_16, s138_17, s138_18, s138_19, s138_20, s138_21, s138_22, s140, s142)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s140, const00000) = '1' then s143_0 <= s142; else s143_0 <= s138_0; end if;
     if equal(s140, const00001) = '1' then s143_1 <= s142; else s143_1 <= s138_1; end if;
     if equal(s140, const00010) = '1' then s143_2 <= s142; else s143_2 <= s138_2; end if;
     if equal(s140, const00011) = '1' then s143_3 <= s142; else s143_3 <= s138_3; end if;
     if equal(s140, const00100) = '1' then s143_4 <= s142; else s143_4 <= s138_4; end if;
     if equal(s140, const00101) = '1' then s143_5 <= s142; else s143_5 <= s138_5; end if;
     if equal(s140, const00110) = '1' then s143_6 <= s142; else s143_6 <= s138_6; end if;
     if equal(s140, const00111) = '1' then s143_7 <= s142; else s143_7 <= s138_7; end if;
     if equal(s140, const01000) = '1' then s143_8 <= s142; else s143_8 <= s138_8; end if;
     if equal(s140, const01001) = '1' then s143_9 <= s142; else s143_9 <= s138_9; end if;
     if equal(s140, const01010) = '1' then s143_10 <= s142; else s143_10 <= s138_10; end if;
     if equal(s140, const01011) = '1' then s143_11 <= s142; else s143_11 <= s138_11; end if;
     if equal(s140, const01100) = '1' then s143_12 <= s142; else s143_12 <= s138_12; end if;
     if equal(s140, const01101) = '1' then s143_13 <= s142; else s143_13 <= s138_13; end if;
     if equal(s140, const01110) = '1' then s143_14 <= s142; else s143_14 <= s138_14; end if;
     if equal(s140, const01111) = '1' then s143_15 <= s142; else s143_15 <= s138_15; end if;
     if equal(s140, const10000) = '1' then s143_16 <= s142; else s143_16 <= s138_16; end if;
     if equal(s140, const10001) = '1' then s143_17 <= s142; else s143_17 <= s138_17; end if;
     if equal(s140, const10010) = '1' then s143_18 <= s142; else s143_18 <= s138_18; end if;
     if equal(s140, const10011) = '1' then s143_19 <= s142; else s143_19 <= s138_19; end if;
     if equal(s140, const10100) = '1' then s143_20 <= s142; else s143_20 <= s138_20; end if;
     if equal(s140, const10101) = '1' then s143_21 <= s142; else s143_21 <= s138_21; end if;
     if equal(s140, const10110) = '1' then s143_22 <= s142; else s143_22 <= s138_22; end if;
   end process;

   s145 <= "00010";  -- constint module constint_2_121

   -- array reader array_reader_122
   process(s143_0, s143_1, s143_2, s143_3, s143_4, s143_5, s143_6, s143_7, s143_8, s143_9, s143_10, s143_11, s143_12, s143_13, s143_14, s143_15, s143_16, s143_17, s143_18, s143_19, s143_20, s143_21, s143_22, s145)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s145, const00000) = '1' ) then s146 <= s143_0; else
       if (equal(s145, const00001) = '1' ) then s146 <= s143_1; else
       if (equal(s145, const00010) = '1' ) then s146 <= s143_2; else
       if (equal(s145, const00011) = '1' ) then s146 <= s143_3; else
       if (equal(s145, const00100) = '1' ) then s146 <= s143_4; else
       if (equal(s145, const00101) = '1' ) then s146 <= s143_5; else
       if (equal(s145, const00110) = '1' ) then s146 <= s143_6; else
       if (equal(s145, const00111) = '1' ) then s146 <= s143_7; else
       if (equal(s145, const01000) = '1' ) then s146 <= s143_8; else
       if (equal(s145, const01001) = '1' ) then s146 <= s143_9; else
       if (equal(s145, const01010) = '1' ) then s146 <= s143_10; else
       if (equal(s145, const01011) = '1' ) then s146 <= s143_11; else
       if (equal(s145, const01100) = '1' ) then s146 <= s143_12; else
       if (equal(s145, const01101) = '1' ) then s146 <= s143_13; else
       if (equal(s145, const01110) = '1' ) then s146 <= s143_14; else
       if (equal(s145, const01111) = '1' ) then s146 <= s143_15; else
       if (equal(s145, const10000) = '1' ) then s146 <= s143_16; else
       if (equal(s145, const10001) = '1' ) then s146 <= s143_17; else
       if (equal(s145, const10010) = '1' ) then s146 <= s143_18; else
       if (equal(s145, const10011) = '1' ) then s146 <= s143_19; else
       if (equal(s145, const10100) = '1' ) then s146 <= s143_20; else
       if (equal(s145, const10101) = '1' ) then s146 <= s143_21; else
       s146 <= s143_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_123
   process(s133, s146, s144)
   begin
   if ( s133 = '1') then s147 <= s144; else s147 <= s146;
   end if;
   end process;

   -- array writer array_writer_124
   process(s143_0, s143_1, s143_2, s143_3, s143_4, s143_5, s143_6, s143_7, s143_8, s143_9, s143_10, s143_11, s143_12, s143_13, s143_14, s143_15, s143_16, s143_17, s143_18, s143_19, s143_20, s143_21, s143_22, s145, s147)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s145, const00000) = '1' then s148_0 <= s147; else s148_0 <= s143_0; end if;
     if equal(s145, const00001) = '1' then s148_1 <= s147; else s148_1 <= s143_1; end if;
     if equal(s145, const00010) = '1' then s148_2 <= s147; else s148_2 <= s143_2; end if;
     if equal(s145, const00011) = '1' then s148_3 <= s147; else s148_3 <= s143_3; end if;
     if equal(s145, const00100) = '1' then s148_4 <= s147; else s148_4 <= s143_4; end if;
     if equal(s145, const00101) = '1' then s148_5 <= s147; else s148_5 <= s143_5; end if;
     if equal(s145, const00110) = '1' then s148_6 <= s147; else s148_6 <= s143_6; end if;
     if equal(s145, const00111) = '1' then s148_7 <= s147; else s148_7 <= s143_7; end if;
     if equal(s145, const01000) = '1' then s148_8 <= s147; else s148_8 <= s143_8; end if;
     if equal(s145, const01001) = '1' then s148_9 <= s147; else s148_9 <= s143_9; end if;
     if equal(s145, const01010) = '1' then s148_10 <= s147; else s148_10 <= s143_10; end if;
     if equal(s145, const01011) = '1' then s148_11 <= s147; else s148_11 <= s143_11; end if;
     if equal(s145, const01100) = '1' then s148_12 <= s147; else s148_12 <= s143_12; end if;
     if equal(s145, const01101) = '1' then s148_13 <= s147; else s148_13 <= s143_13; end if;
     if equal(s145, const01110) = '1' then s148_14 <= s147; else s148_14 <= s143_14; end if;
     if equal(s145, const01111) = '1' then s148_15 <= s147; else s148_15 <= s143_15; end if;
     if equal(s145, const10000) = '1' then s148_16 <= s147; else s148_16 <= s143_16; end if;
     if equal(s145, const10001) = '1' then s148_17 <= s147; else s148_17 <= s143_17; end if;
     if equal(s145, const10010) = '1' then s148_18 <= s147; else s148_18 <= s143_18; end if;
     if equal(s145, const10011) = '1' then s148_19 <= s147; else s148_19 <= s143_19; end if;
     if equal(s145, const10100) = '1' then s148_20 <= s147; else s148_20 <= s143_20; end if;
     if equal(s145, const10101) = '1' then s148_21 <= s147; else s148_21 <= s143_21; end if;
     if equal(s145, const10110) = '1' then s148_22 <= s147; else s148_22 <= s143_22; end if;
   end process;

   s150 <= "00011";  -- constint module constint_3_125

   -- array reader array_reader_126
   process(s148_0, s148_1, s148_2, s148_3, s148_4, s148_5, s148_6, s148_7, s148_8, s148_9, s148_10, s148_11, s148_12, s148_13, s148_14, s148_15, s148_16, s148_17, s148_18, s148_19, s148_20, s148_21, s148_22, s150)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s150, const00000) = '1' ) then s151 <= s148_0; else
       if (equal(s150, const00001) = '1' ) then s151 <= s148_1; else
       if (equal(s150, const00010) = '1' ) then s151 <= s148_2; else
       if (equal(s150, const00011) = '1' ) then s151 <= s148_3; else
       if (equal(s150, const00100) = '1' ) then s151 <= s148_4; else
       if (equal(s150, const00101) = '1' ) then s151 <= s148_5; else
       if (equal(s150, const00110) = '1' ) then s151 <= s148_6; else
       if (equal(s150, const00111) = '1' ) then s151 <= s148_7; else
       if (equal(s150, const01000) = '1' ) then s151 <= s148_8; else
       if (equal(s150, const01001) = '1' ) then s151 <= s148_9; else
       if (equal(s150, const01010) = '1' ) then s151 <= s148_10; else
       if (equal(s150, const01011) = '1' ) then s151 <= s148_11; else
       if (equal(s150, const01100) = '1' ) then s151 <= s148_12; else
       if (equal(s150, const01101) = '1' ) then s151 <= s148_13; else
       if (equal(s150, const01110) = '1' ) then s151 <= s148_14; else
       if (equal(s150, const01111) = '1' ) then s151 <= s148_15; else
       if (equal(s150, const10000) = '1' ) then s151 <= s148_16; else
       if (equal(s150, const10001) = '1' ) then s151 <= s148_17; else
       if (equal(s150, const10010) = '1' ) then s151 <= s148_18; else
       if (equal(s150, const10011) = '1' ) then s151 <= s148_19; else
       if (equal(s150, const10100) = '1' ) then s151 <= s148_20; else
       if (equal(s150, const10101) = '1' ) then s151 <= s148_21; else
       s151 <= s148_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_127
   process(s133, s151, s149)
   begin
   if ( s133 = '1') then s152 <= s149; else s152 <= s151;
   end if;
   end process;

   -- array writer array_writer_128
   process(s148_0, s148_1, s148_2, s148_3, s148_4, s148_5, s148_6, s148_7, s148_8, s148_9, s148_10, s148_11, s148_12, s148_13, s148_14, s148_15, s148_16, s148_17, s148_18, s148_19, s148_20, s148_21, s148_22, s150, s152)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s150, const00000) = '1' then s153_0 <= s152; else s153_0 <= s148_0; end if;
     if equal(s150, const00001) = '1' then s153_1 <= s152; else s153_1 <= s148_1; end if;
     if equal(s150, const00010) = '1' then s153_2 <= s152; else s153_2 <= s148_2; end if;
     if equal(s150, const00011) = '1' then s153_3 <= s152; else s153_3 <= s148_3; end if;
     if equal(s150, const00100) = '1' then s153_4 <= s152; else s153_4 <= s148_4; end if;
     if equal(s150, const00101) = '1' then s153_5 <= s152; else s153_5 <= s148_5; end if;
     if equal(s150, const00110) = '1' then s153_6 <= s152; else s153_6 <= s148_6; end if;
     if equal(s150, const00111) = '1' then s153_7 <= s152; else s153_7 <= s148_7; end if;
     if equal(s150, const01000) = '1' then s153_8 <= s152; else s153_8 <= s148_8; end if;
     if equal(s150, const01001) = '1' then s153_9 <= s152; else s153_9 <= s148_9; end if;
     if equal(s150, const01010) = '1' then s153_10 <= s152; else s153_10 <= s148_10; end if;
     if equal(s150, const01011) = '1' then s153_11 <= s152; else s153_11 <= s148_11; end if;
     if equal(s150, const01100) = '1' then s153_12 <= s152; else s153_12 <= s148_12; end if;
     if equal(s150, const01101) = '1' then s153_13 <= s152; else s153_13 <= s148_13; end if;
     if equal(s150, const01110) = '1' then s153_14 <= s152; else s153_14 <= s148_14; end if;
     if equal(s150, const01111) = '1' then s153_15 <= s152; else s153_15 <= s148_15; end if;
     if equal(s150, const10000) = '1' then s153_16 <= s152; else s153_16 <= s148_16; end if;
     if equal(s150, const10001) = '1' then s153_17 <= s152; else s153_17 <= s148_17; end if;
     if equal(s150, const10010) = '1' then s153_18 <= s152; else s153_18 <= s148_18; end if;
     if equal(s150, const10011) = '1' then s153_19 <= s152; else s153_19 <= s148_19; end if;
     if equal(s150, const10100) = '1' then s153_20 <= s152; else s153_20 <= s148_20; end if;
     if equal(s150, const10101) = '1' then s153_21 <= s152; else s153_21 <= s148_21; end if;
     if equal(s150, const10110) = '1' then s153_22 <= s152; else s153_22 <= s148_22; end if;
   end process;

   s155 <= "00100";  -- constint module constint_4_129

   -- array reader array_reader_130
   process(s153_0, s153_1, s153_2, s153_3, s153_4, s153_5, s153_6, s153_7, s153_8, s153_9, s153_10, s153_11, s153_12, s153_13, s153_14, s153_15, s153_16, s153_17, s153_18, s153_19, s153_20, s153_21, s153_22, s155)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s155, const00000) = '1' ) then s156 <= s153_0; else
       if (equal(s155, const00001) = '1' ) then s156 <= s153_1; else
       if (equal(s155, const00010) = '1' ) then s156 <= s153_2; else
       if (equal(s155, const00011) = '1' ) then s156 <= s153_3; else
       if (equal(s155, const00100) = '1' ) then s156 <= s153_4; else
       if (equal(s155, const00101) = '1' ) then s156 <= s153_5; else
       if (equal(s155, const00110) = '1' ) then s156 <= s153_6; else
       if (equal(s155, const00111) = '1' ) then s156 <= s153_7; else
       if (equal(s155, const01000) = '1' ) then s156 <= s153_8; else
       if (equal(s155, const01001) = '1' ) then s156 <= s153_9; else
       if (equal(s155, const01010) = '1' ) then s156 <= s153_10; else
       if (equal(s155, const01011) = '1' ) then s156 <= s153_11; else
       if (equal(s155, const01100) = '1' ) then s156 <= s153_12; else
       if (equal(s155, const01101) = '1' ) then s156 <= s153_13; else
       if (equal(s155, const01110) = '1' ) then s156 <= s153_14; else
       if (equal(s155, const01111) = '1' ) then s156 <= s153_15; else
       if (equal(s155, const10000) = '1' ) then s156 <= s153_16; else
       if (equal(s155, const10001) = '1' ) then s156 <= s153_17; else
       if (equal(s155, const10010) = '1' ) then s156 <= s153_18; else
       if (equal(s155, const10011) = '1' ) then s156 <= s153_19; else
       if (equal(s155, const10100) = '1' ) then s156 <= s153_20; else
       if (equal(s155, const10101) = '1' ) then s156 <= s153_21; else
       s156 <= s153_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_131
   process(s133, s156, s154)
   begin
   if ( s133 = '1') then s157 <= s154; else s157 <= s156;
   end if;
   end process;

   -- array writer array_writer_132
   process(s153_0, s153_1, s153_2, s153_3, s153_4, s153_5, s153_6, s153_7, s153_8, s153_9, s153_10, s153_11, s153_12, s153_13, s153_14, s153_15, s153_16, s153_17, s153_18, s153_19, s153_20, s153_21, s153_22, s155, s157)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s155, const00000) = '1' then s158_0 <= s157; else s158_0 <= s153_0; end if;
     if equal(s155, const00001) = '1' then s158_1 <= s157; else s158_1 <= s153_1; end if;
     if equal(s155, const00010) = '1' then s158_2 <= s157; else s158_2 <= s153_2; end if;
     if equal(s155, const00011) = '1' then s158_3 <= s157; else s158_3 <= s153_3; end if;
     if equal(s155, const00100) = '1' then s158_4 <= s157; else s158_4 <= s153_4; end if;
     if equal(s155, const00101) = '1' then s158_5 <= s157; else s158_5 <= s153_5; end if;
     if equal(s155, const00110) = '1' then s158_6 <= s157; else s158_6 <= s153_6; end if;
     if equal(s155, const00111) = '1' then s158_7 <= s157; else s158_7 <= s153_7; end if;
     if equal(s155, const01000) = '1' then s158_8 <= s157; else s158_8 <= s153_8; end if;
     if equal(s155, const01001) = '1' then s158_9 <= s157; else s158_9 <= s153_9; end if;
     if equal(s155, const01010) = '1' then s158_10 <= s157; else s158_10 <= s153_10; end if;
     if equal(s155, const01011) = '1' then s158_11 <= s157; else s158_11 <= s153_11; end if;
     if equal(s155, const01100) = '1' then s158_12 <= s157; else s158_12 <= s153_12; end if;
     if equal(s155, const01101) = '1' then s158_13 <= s157; else s158_13 <= s153_13; end if;
     if equal(s155, const01110) = '1' then s158_14 <= s157; else s158_14 <= s153_14; end if;
     if equal(s155, const01111) = '1' then s158_15 <= s157; else s158_15 <= s153_15; end if;
     if equal(s155, const10000) = '1' then s158_16 <= s157; else s158_16 <= s153_16; end if;
     if equal(s155, const10001) = '1' then s158_17 <= s157; else s158_17 <= s153_17; end if;
     if equal(s155, const10010) = '1' then s158_18 <= s157; else s158_18 <= s153_18; end if;
     if equal(s155, const10011) = '1' then s158_19 <= s157; else s158_19 <= s153_19; end if;
     if equal(s155, const10100) = '1' then s158_20 <= s157; else s158_20 <= s153_20; end if;
     if equal(s155, const10101) = '1' then s158_21 <= s157; else s158_21 <= s153_21; end if;
     if equal(s155, const10110) = '1' then s158_22 <= s157; else s158_22 <= s153_22; end if;
   end process;

   s160 <= "00101";  -- constint module constint_5_133

   -- array reader array_reader_134
   process(s158_0, s158_1, s158_2, s158_3, s158_4, s158_5, s158_6, s158_7, s158_8, s158_9, s158_10, s158_11, s158_12, s158_13, s158_14, s158_15, s158_16, s158_17, s158_18, s158_19, s158_20, s158_21, s158_22, s160)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s160, const00000) = '1' ) then s161 <= s158_0; else
       if (equal(s160, const00001) = '1' ) then s161 <= s158_1; else
       if (equal(s160, const00010) = '1' ) then s161 <= s158_2; else
       if (equal(s160, const00011) = '1' ) then s161 <= s158_3; else
       if (equal(s160, const00100) = '1' ) then s161 <= s158_4; else
       if (equal(s160, const00101) = '1' ) then s161 <= s158_5; else
       if (equal(s160, const00110) = '1' ) then s161 <= s158_6; else
       if (equal(s160, const00111) = '1' ) then s161 <= s158_7; else
       if (equal(s160, const01000) = '1' ) then s161 <= s158_8; else
       if (equal(s160, const01001) = '1' ) then s161 <= s158_9; else
       if (equal(s160, const01010) = '1' ) then s161 <= s158_10; else
       if (equal(s160, const01011) = '1' ) then s161 <= s158_11; else
       if (equal(s160, const01100) = '1' ) then s161 <= s158_12; else
       if (equal(s160, const01101) = '1' ) then s161 <= s158_13; else
       if (equal(s160, const01110) = '1' ) then s161 <= s158_14; else
       if (equal(s160, const01111) = '1' ) then s161 <= s158_15; else
       if (equal(s160, const10000) = '1' ) then s161 <= s158_16; else
       if (equal(s160, const10001) = '1' ) then s161 <= s158_17; else
       if (equal(s160, const10010) = '1' ) then s161 <= s158_18; else
       if (equal(s160, const10011) = '1' ) then s161 <= s158_19; else
       if (equal(s160, const10100) = '1' ) then s161 <= s158_20; else
       if (equal(s160, const10101) = '1' ) then s161 <= s158_21; else
       s161 <= s158_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_135
   process(s133, s161, s159)
   begin
   if ( s133 = '1') then s162 <= s159; else s162 <= s161;
   end if;
   end process;

   -- array writer array_writer_136
   process(s158_0, s158_1, s158_2, s158_3, s158_4, s158_5, s158_6, s158_7, s158_8, s158_9, s158_10, s158_11, s158_12, s158_13, s158_14, s158_15, s158_16, s158_17, s158_18, s158_19, s158_20, s158_21, s158_22, s160, s162)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s160, const00000) = '1' then s163_0 <= s162; else s163_0 <= s158_0; end if;
     if equal(s160, const00001) = '1' then s163_1 <= s162; else s163_1 <= s158_1; end if;
     if equal(s160, const00010) = '1' then s163_2 <= s162; else s163_2 <= s158_2; end if;
     if equal(s160, const00011) = '1' then s163_3 <= s162; else s163_3 <= s158_3; end if;
     if equal(s160, const00100) = '1' then s163_4 <= s162; else s163_4 <= s158_4; end if;
     if equal(s160, const00101) = '1' then s163_5 <= s162; else s163_5 <= s158_5; end if;
     if equal(s160, const00110) = '1' then s163_6 <= s162; else s163_6 <= s158_6; end if;
     if equal(s160, const00111) = '1' then s163_7 <= s162; else s163_7 <= s158_7; end if;
     if equal(s160, const01000) = '1' then s163_8 <= s162; else s163_8 <= s158_8; end if;
     if equal(s160, const01001) = '1' then s163_9 <= s162; else s163_9 <= s158_9; end if;
     if equal(s160, const01010) = '1' then s163_10 <= s162; else s163_10 <= s158_10; end if;
     if equal(s160, const01011) = '1' then s163_11 <= s162; else s163_11 <= s158_11; end if;
     if equal(s160, const01100) = '1' then s163_12 <= s162; else s163_12 <= s158_12; end if;
     if equal(s160, const01101) = '1' then s163_13 <= s162; else s163_13 <= s158_13; end if;
     if equal(s160, const01110) = '1' then s163_14 <= s162; else s163_14 <= s158_14; end if;
     if equal(s160, const01111) = '1' then s163_15 <= s162; else s163_15 <= s158_15; end if;
     if equal(s160, const10000) = '1' then s163_16 <= s162; else s163_16 <= s158_16; end if;
     if equal(s160, const10001) = '1' then s163_17 <= s162; else s163_17 <= s158_17; end if;
     if equal(s160, const10010) = '1' then s163_18 <= s162; else s163_18 <= s158_18; end if;
     if equal(s160, const10011) = '1' then s163_19 <= s162; else s163_19 <= s158_19; end if;
     if equal(s160, const10100) = '1' then s163_20 <= s162; else s163_20 <= s158_20; end if;
     if equal(s160, const10101) = '1' then s163_21 <= s162; else s163_21 <= s158_21; end if;
     if equal(s160, const10110) = '1' then s163_22 <= s162; else s163_22 <= s158_22; end if;
   end process;

   s165 <= "00110";  -- constint module constint_6_137

   -- array reader array_reader_138
   process(s163_0, s163_1, s163_2, s163_3, s163_4, s163_5, s163_6, s163_7, s163_8, s163_9, s163_10, s163_11, s163_12, s163_13, s163_14, s163_15, s163_16, s163_17, s163_18, s163_19, s163_20, s163_21, s163_22, s165)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s165, const00000) = '1' ) then s166 <= s163_0; else
       if (equal(s165, const00001) = '1' ) then s166 <= s163_1; else
       if (equal(s165, const00010) = '1' ) then s166 <= s163_2; else
       if (equal(s165, const00011) = '1' ) then s166 <= s163_3; else
       if (equal(s165, const00100) = '1' ) then s166 <= s163_4; else
       if (equal(s165, const00101) = '1' ) then s166 <= s163_5; else
       if (equal(s165, const00110) = '1' ) then s166 <= s163_6; else
       if (equal(s165, const00111) = '1' ) then s166 <= s163_7; else
       if (equal(s165, const01000) = '1' ) then s166 <= s163_8; else
       if (equal(s165, const01001) = '1' ) then s166 <= s163_9; else
       if (equal(s165, const01010) = '1' ) then s166 <= s163_10; else
       if (equal(s165, const01011) = '1' ) then s166 <= s163_11; else
       if (equal(s165, const01100) = '1' ) then s166 <= s163_12; else
       if (equal(s165, const01101) = '1' ) then s166 <= s163_13; else
       if (equal(s165, const01110) = '1' ) then s166 <= s163_14; else
       if (equal(s165, const01111) = '1' ) then s166 <= s163_15; else
       if (equal(s165, const10000) = '1' ) then s166 <= s163_16; else
       if (equal(s165, const10001) = '1' ) then s166 <= s163_17; else
       if (equal(s165, const10010) = '1' ) then s166 <= s163_18; else
       if (equal(s165, const10011) = '1' ) then s166 <= s163_19; else
       if (equal(s165, const10100) = '1' ) then s166 <= s163_20; else
       if (equal(s165, const10101) = '1' ) then s166 <= s163_21; else
       s166 <= s163_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_139
   process(s133, s166, s164)
   begin
   if ( s133 = '1') then s167 <= s164; else s167 <= s166;
   end if;
   end process;

   -- array writer array_writer_140
   process(s163_0, s163_1, s163_2, s163_3, s163_4, s163_5, s163_6, s163_7, s163_8, s163_9, s163_10, s163_11, s163_12, s163_13, s163_14, s163_15, s163_16, s163_17, s163_18, s163_19, s163_20, s163_21, s163_22, s165, s167)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s165, const00000) = '1' then s168_0 <= s167; else s168_0 <= s163_0; end if;
     if equal(s165, const00001) = '1' then s168_1 <= s167; else s168_1 <= s163_1; end if;
     if equal(s165, const00010) = '1' then s168_2 <= s167; else s168_2 <= s163_2; end if;
     if equal(s165, const00011) = '1' then s168_3 <= s167; else s168_3 <= s163_3; end if;
     if equal(s165, const00100) = '1' then s168_4 <= s167; else s168_4 <= s163_4; end if;
     if equal(s165, const00101) = '1' then s168_5 <= s167; else s168_5 <= s163_5; end if;
     if equal(s165, const00110) = '1' then s168_6 <= s167; else s168_6 <= s163_6; end if;
     if equal(s165, const00111) = '1' then s168_7 <= s167; else s168_7 <= s163_7; end if;
     if equal(s165, const01000) = '1' then s168_8 <= s167; else s168_8 <= s163_8; end if;
     if equal(s165, const01001) = '1' then s168_9 <= s167; else s168_9 <= s163_9; end if;
     if equal(s165, const01010) = '1' then s168_10 <= s167; else s168_10 <= s163_10; end if;
     if equal(s165, const01011) = '1' then s168_11 <= s167; else s168_11 <= s163_11; end if;
     if equal(s165, const01100) = '1' then s168_12 <= s167; else s168_12 <= s163_12; end if;
     if equal(s165, const01101) = '1' then s168_13 <= s167; else s168_13 <= s163_13; end if;
     if equal(s165, const01110) = '1' then s168_14 <= s167; else s168_14 <= s163_14; end if;
     if equal(s165, const01111) = '1' then s168_15 <= s167; else s168_15 <= s163_15; end if;
     if equal(s165, const10000) = '1' then s168_16 <= s167; else s168_16 <= s163_16; end if;
     if equal(s165, const10001) = '1' then s168_17 <= s167; else s168_17 <= s163_17; end if;
     if equal(s165, const10010) = '1' then s168_18 <= s167; else s168_18 <= s163_18; end if;
     if equal(s165, const10011) = '1' then s168_19 <= s167; else s168_19 <= s163_19; end if;
     if equal(s165, const10100) = '1' then s168_20 <= s167; else s168_20 <= s163_20; end if;
     if equal(s165, const10101) = '1' then s168_21 <= s167; else s168_21 <= s163_21; end if;
     if equal(s165, const10110) = '1' then s168_22 <= s167; else s168_22 <= s163_22; end if;
   end process;

   s170 <= "00111";  -- constint module constint_7_141

   -- array reader array_reader_142
   process(s168_0, s168_1, s168_2, s168_3, s168_4, s168_5, s168_6, s168_7, s168_8, s168_9, s168_10, s168_11, s168_12, s168_13, s168_14, s168_15, s168_16, s168_17, s168_18, s168_19, s168_20, s168_21, s168_22, s170)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s170, const00000) = '1' ) then s171 <= s168_0; else
       if (equal(s170, const00001) = '1' ) then s171 <= s168_1; else
       if (equal(s170, const00010) = '1' ) then s171 <= s168_2; else
       if (equal(s170, const00011) = '1' ) then s171 <= s168_3; else
       if (equal(s170, const00100) = '1' ) then s171 <= s168_4; else
       if (equal(s170, const00101) = '1' ) then s171 <= s168_5; else
       if (equal(s170, const00110) = '1' ) then s171 <= s168_6; else
       if (equal(s170, const00111) = '1' ) then s171 <= s168_7; else
       if (equal(s170, const01000) = '1' ) then s171 <= s168_8; else
       if (equal(s170, const01001) = '1' ) then s171 <= s168_9; else
       if (equal(s170, const01010) = '1' ) then s171 <= s168_10; else
       if (equal(s170, const01011) = '1' ) then s171 <= s168_11; else
       if (equal(s170, const01100) = '1' ) then s171 <= s168_12; else
       if (equal(s170, const01101) = '1' ) then s171 <= s168_13; else
       if (equal(s170, const01110) = '1' ) then s171 <= s168_14; else
       if (equal(s170, const01111) = '1' ) then s171 <= s168_15; else
       if (equal(s170, const10000) = '1' ) then s171 <= s168_16; else
       if (equal(s170, const10001) = '1' ) then s171 <= s168_17; else
       if (equal(s170, const10010) = '1' ) then s171 <= s168_18; else
       if (equal(s170, const10011) = '1' ) then s171 <= s168_19; else
       if (equal(s170, const10100) = '1' ) then s171 <= s168_20; else
       if (equal(s170, const10101) = '1' ) then s171 <= s168_21; else
       s171 <= s168_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_143
   process(s133, s171, s169)
   begin
   if ( s133 = '1') then s172 <= s169; else s172 <= s171;
   end if;
   end process;

   -- array writer array_writer_144
   process(s168_0, s168_1, s168_2, s168_3, s168_4, s168_5, s168_6, s168_7, s168_8, s168_9, s168_10, s168_11, s168_12, s168_13, s168_14, s168_15, s168_16, s168_17, s168_18, s168_19, s168_20, s168_21, s168_22, s170, s172)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s170, const00000) = '1' then s173_0 <= s172; else s173_0 <= s168_0; end if;
     if equal(s170, const00001) = '1' then s173_1 <= s172; else s173_1 <= s168_1; end if;
     if equal(s170, const00010) = '1' then s173_2 <= s172; else s173_2 <= s168_2; end if;
     if equal(s170, const00011) = '1' then s173_3 <= s172; else s173_3 <= s168_3; end if;
     if equal(s170, const00100) = '1' then s173_4 <= s172; else s173_4 <= s168_4; end if;
     if equal(s170, const00101) = '1' then s173_5 <= s172; else s173_5 <= s168_5; end if;
     if equal(s170, const00110) = '1' then s173_6 <= s172; else s173_6 <= s168_6; end if;
     if equal(s170, const00111) = '1' then s173_7 <= s172; else s173_7 <= s168_7; end if;
     if equal(s170, const01000) = '1' then s173_8 <= s172; else s173_8 <= s168_8; end if;
     if equal(s170, const01001) = '1' then s173_9 <= s172; else s173_9 <= s168_9; end if;
     if equal(s170, const01010) = '1' then s173_10 <= s172; else s173_10 <= s168_10; end if;
     if equal(s170, const01011) = '1' then s173_11 <= s172; else s173_11 <= s168_11; end if;
     if equal(s170, const01100) = '1' then s173_12 <= s172; else s173_12 <= s168_12; end if;
     if equal(s170, const01101) = '1' then s173_13 <= s172; else s173_13 <= s168_13; end if;
     if equal(s170, const01110) = '1' then s173_14 <= s172; else s173_14 <= s168_14; end if;
     if equal(s170, const01111) = '1' then s173_15 <= s172; else s173_15 <= s168_15; end if;
     if equal(s170, const10000) = '1' then s173_16 <= s172; else s173_16 <= s168_16; end if;
     if equal(s170, const10001) = '1' then s173_17 <= s172; else s173_17 <= s168_17; end if;
     if equal(s170, const10010) = '1' then s173_18 <= s172; else s173_18 <= s168_18; end if;
     if equal(s170, const10011) = '1' then s173_19 <= s172; else s173_19 <= s168_19; end if;
     if equal(s170, const10100) = '1' then s173_20 <= s172; else s173_20 <= s168_20; end if;
     if equal(s170, const10101) = '1' then s173_21 <= s172; else s173_21 <= s168_21; end if;
     if equal(s170, const10110) = '1' then s173_22 <= s172; else s173_22 <= s168_22; end if;
   end process;

   s175 <= "01000";  -- constint module constint_8_145

   -- array reader array_reader_146
   process(s173_0, s173_1, s173_2, s173_3, s173_4, s173_5, s173_6, s173_7, s173_8, s173_9, s173_10, s173_11, s173_12, s173_13, s173_14, s173_15, s173_16, s173_17, s173_18, s173_19, s173_20, s173_21, s173_22, s175)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s175, const00000) = '1' ) then s176 <= s173_0; else
       if (equal(s175, const00001) = '1' ) then s176 <= s173_1; else
       if (equal(s175, const00010) = '1' ) then s176 <= s173_2; else
       if (equal(s175, const00011) = '1' ) then s176 <= s173_3; else
       if (equal(s175, const00100) = '1' ) then s176 <= s173_4; else
       if (equal(s175, const00101) = '1' ) then s176 <= s173_5; else
       if (equal(s175, const00110) = '1' ) then s176 <= s173_6; else
       if (equal(s175, const00111) = '1' ) then s176 <= s173_7; else
       if (equal(s175, const01000) = '1' ) then s176 <= s173_8; else
       if (equal(s175, const01001) = '1' ) then s176 <= s173_9; else
       if (equal(s175, const01010) = '1' ) then s176 <= s173_10; else
       if (equal(s175, const01011) = '1' ) then s176 <= s173_11; else
       if (equal(s175, const01100) = '1' ) then s176 <= s173_12; else
       if (equal(s175, const01101) = '1' ) then s176 <= s173_13; else
       if (equal(s175, const01110) = '1' ) then s176 <= s173_14; else
       if (equal(s175, const01111) = '1' ) then s176 <= s173_15; else
       if (equal(s175, const10000) = '1' ) then s176 <= s173_16; else
       if (equal(s175, const10001) = '1' ) then s176 <= s173_17; else
       if (equal(s175, const10010) = '1' ) then s176 <= s173_18; else
       if (equal(s175, const10011) = '1' ) then s176 <= s173_19; else
       if (equal(s175, const10100) = '1' ) then s176 <= s173_20; else
       if (equal(s175, const10101) = '1' ) then s176 <= s173_21; else
       s176 <= s173_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_147
   process(s133, s176, s174)
   begin
   if ( s133 = '1') then s177 <= s174; else s177 <= s176;
   end if;
   end process;

   -- array writer array_writer_148
   process(s173_0, s173_1, s173_2, s173_3, s173_4, s173_5, s173_6, s173_7, s173_8, s173_9, s173_10, s173_11, s173_12, s173_13, s173_14, s173_15, s173_16, s173_17, s173_18, s173_19, s173_20, s173_21, s173_22, s175, s177)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s175, const00000) = '1' then s178_0 <= s177; else s178_0 <= s173_0; end if;
     if equal(s175, const00001) = '1' then s178_1 <= s177; else s178_1 <= s173_1; end if;
     if equal(s175, const00010) = '1' then s178_2 <= s177; else s178_2 <= s173_2; end if;
     if equal(s175, const00011) = '1' then s178_3 <= s177; else s178_3 <= s173_3; end if;
     if equal(s175, const00100) = '1' then s178_4 <= s177; else s178_4 <= s173_4; end if;
     if equal(s175, const00101) = '1' then s178_5 <= s177; else s178_5 <= s173_5; end if;
     if equal(s175, const00110) = '1' then s178_6 <= s177; else s178_6 <= s173_6; end if;
     if equal(s175, const00111) = '1' then s178_7 <= s177; else s178_7 <= s173_7; end if;
     if equal(s175, const01000) = '1' then s178_8 <= s177; else s178_8 <= s173_8; end if;
     if equal(s175, const01001) = '1' then s178_9 <= s177; else s178_9 <= s173_9; end if;
     if equal(s175, const01010) = '1' then s178_10 <= s177; else s178_10 <= s173_10; end if;
     if equal(s175, const01011) = '1' then s178_11 <= s177; else s178_11 <= s173_11; end if;
     if equal(s175, const01100) = '1' then s178_12 <= s177; else s178_12 <= s173_12; end if;
     if equal(s175, const01101) = '1' then s178_13 <= s177; else s178_13 <= s173_13; end if;
     if equal(s175, const01110) = '1' then s178_14 <= s177; else s178_14 <= s173_14; end if;
     if equal(s175, const01111) = '1' then s178_15 <= s177; else s178_15 <= s173_15; end if;
     if equal(s175, const10000) = '1' then s178_16 <= s177; else s178_16 <= s173_16; end if;
     if equal(s175, const10001) = '1' then s178_17 <= s177; else s178_17 <= s173_17; end if;
     if equal(s175, const10010) = '1' then s178_18 <= s177; else s178_18 <= s173_18; end if;
     if equal(s175, const10011) = '1' then s178_19 <= s177; else s178_19 <= s173_19; end if;
     if equal(s175, const10100) = '1' then s178_20 <= s177; else s178_20 <= s173_20; end if;
     if equal(s175, const10101) = '1' then s178_21 <= s177; else s178_21 <= s173_21; end if;
     if equal(s175, const10110) = '1' then s178_22 <= s177; else s178_22 <= s173_22; end if;
   end process;

   s180 <= "01001";  -- constint module constint_9_149

   -- array reader array_reader_150
   process(s178_0, s178_1, s178_2, s178_3, s178_4, s178_5, s178_6, s178_7, s178_8, s178_9, s178_10, s178_11, s178_12, s178_13, s178_14, s178_15, s178_16, s178_17, s178_18, s178_19, s178_20, s178_21, s178_22, s180)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s180, const00000) = '1' ) then s181 <= s178_0; else
       if (equal(s180, const00001) = '1' ) then s181 <= s178_1; else
       if (equal(s180, const00010) = '1' ) then s181 <= s178_2; else
       if (equal(s180, const00011) = '1' ) then s181 <= s178_3; else
       if (equal(s180, const00100) = '1' ) then s181 <= s178_4; else
       if (equal(s180, const00101) = '1' ) then s181 <= s178_5; else
       if (equal(s180, const00110) = '1' ) then s181 <= s178_6; else
       if (equal(s180, const00111) = '1' ) then s181 <= s178_7; else
       if (equal(s180, const01000) = '1' ) then s181 <= s178_8; else
       if (equal(s180, const01001) = '1' ) then s181 <= s178_9; else
       if (equal(s180, const01010) = '1' ) then s181 <= s178_10; else
       if (equal(s180, const01011) = '1' ) then s181 <= s178_11; else
       if (equal(s180, const01100) = '1' ) then s181 <= s178_12; else
       if (equal(s180, const01101) = '1' ) then s181 <= s178_13; else
       if (equal(s180, const01110) = '1' ) then s181 <= s178_14; else
       if (equal(s180, const01111) = '1' ) then s181 <= s178_15; else
       if (equal(s180, const10000) = '1' ) then s181 <= s178_16; else
       if (equal(s180, const10001) = '1' ) then s181 <= s178_17; else
       if (equal(s180, const10010) = '1' ) then s181 <= s178_18; else
       if (equal(s180, const10011) = '1' ) then s181 <= s178_19; else
       if (equal(s180, const10100) = '1' ) then s181 <= s178_20; else
       if (equal(s180, const10101) = '1' ) then s181 <= s178_21; else
       s181 <= s178_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_151
   process(s133, s181, s179)
   begin
   if ( s133 = '1') then s182 <= s179; else s182 <= s181;
   end if;
   end process;

   -- array writer array_writer_152
   process(s178_0, s178_1, s178_2, s178_3, s178_4, s178_5, s178_6, s178_7, s178_8, s178_9, s178_10, s178_11, s178_12, s178_13, s178_14, s178_15, s178_16, s178_17, s178_18, s178_19, s178_20, s178_21, s178_22, s180, s182)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s180, const00000) = '1' then s183_0 <= s182; else s183_0 <= s178_0; end if;
     if equal(s180, const00001) = '1' then s183_1 <= s182; else s183_1 <= s178_1; end if;
     if equal(s180, const00010) = '1' then s183_2 <= s182; else s183_2 <= s178_2; end if;
     if equal(s180, const00011) = '1' then s183_3 <= s182; else s183_3 <= s178_3; end if;
     if equal(s180, const00100) = '1' then s183_4 <= s182; else s183_4 <= s178_4; end if;
     if equal(s180, const00101) = '1' then s183_5 <= s182; else s183_5 <= s178_5; end if;
     if equal(s180, const00110) = '1' then s183_6 <= s182; else s183_6 <= s178_6; end if;
     if equal(s180, const00111) = '1' then s183_7 <= s182; else s183_7 <= s178_7; end if;
     if equal(s180, const01000) = '1' then s183_8 <= s182; else s183_8 <= s178_8; end if;
     if equal(s180, const01001) = '1' then s183_9 <= s182; else s183_9 <= s178_9; end if;
     if equal(s180, const01010) = '1' then s183_10 <= s182; else s183_10 <= s178_10; end if;
     if equal(s180, const01011) = '1' then s183_11 <= s182; else s183_11 <= s178_11; end if;
     if equal(s180, const01100) = '1' then s183_12 <= s182; else s183_12 <= s178_12; end if;
     if equal(s180, const01101) = '1' then s183_13 <= s182; else s183_13 <= s178_13; end if;
     if equal(s180, const01110) = '1' then s183_14 <= s182; else s183_14 <= s178_14; end if;
     if equal(s180, const01111) = '1' then s183_15 <= s182; else s183_15 <= s178_15; end if;
     if equal(s180, const10000) = '1' then s183_16 <= s182; else s183_16 <= s178_16; end if;
     if equal(s180, const10001) = '1' then s183_17 <= s182; else s183_17 <= s178_17; end if;
     if equal(s180, const10010) = '1' then s183_18 <= s182; else s183_18 <= s178_18; end if;
     if equal(s180, const10011) = '1' then s183_19 <= s182; else s183_19 <= s178_19; end if;
     if equal(s180, const10100) = '1' then s183_20 <= s182; else s183_20 <= s178_20; end if;
     if equal(s180, const10101) = '1' then s183_21 <= s182; else s183_21 <= s178_21; end if;
     if equal(s180, const10110) = '1' then s183_22 <= s182; else s183_22 <= s178_22; end if;
   end process;

   s185 <= "01010";  -- constint module constint_10_153

   -- array reader array_reader_154
   process(s183_0, s183_1, s183_2, s183_3, s183_4, s183_5, s183_6, s183_7, s183_8, s183_9, s183_10, s183_11, s183_12, s183_13, s183_14, s183_15, s183_16, s183_17, s183_18, s183_19, s183_20, s183_21, s183_22, s185)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s185, const00000) = '1' ) then s186 <= s183_0; else
       if (equal(s185, const00001) = '1' ) then s186 <= s183_1; else
       if (equal(s185, const00010) = '1' ) then s186 <= s183_2; else
       if (equal(s185, const00011) = '1' ) then s186 <= s183_3; else
       if (equal(s185, const00100) = '1' ) then s186 <= s183_4; else
       if (equal(s185, const00101) = '1' ) then s186 <= s183_5; else
       if (equal(s185, const00110) = '1' ) then s186 <= s183_6; else
       if (equal(s185, const00111) = '1' ) then s186 <= s183_7; else
       if (equal(s185, const01000) = '1' ) then s186 <= s183_8; else
       if (equal(s185, const01001) = '1' ) then s186 <= s183_9; else
       if (equal(s185, const01010) = '1' ) then s186 <= s183_10; else
       if (equal(s185, const01011) = '1' ) then s186 <= s183_11; else
       if (equal(s185, const01100) = '1' ) then s186 <= s183_12; else
       if (equal(s185, const01101) = '1' ) then s186 <= s183_13; else
       if (equal(s185, const01110) = '1' ) then s186 <= s183_14; else
       if (equal(s185, const01111) = '1' ) then s186 <= s183_15; else
       if (equal(s185, const10000) = '1' ) then s186 <= s183_16; else
       if (equal(s185, const10001) = '1' ) then s186 <= s183_17; else
       if (equal(s185, const10010) = '1' ) then s186 <= s183_18; else
       if (equal(s185, const10011) = '1' ) then s186 <= s183_19; else
       if (equal(s185, const10100) = '1' ) then s186 <= s183_20; else
       if (equal(s185, const10101) = '1' ) then s186 <= s183_21; else
       s186 <= s183_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_155
   process(s133, s186, s184)
   begin
   if ( s133 = '1') then s187 <= s184; else s187 <= s186;
   end if;
   end process;

   -- array writer array_writer_156
   process(s183_0, s183_1, s183_2, s183_3, s183_4, s183_5, s183_6, s183_7, s183_8, s183_9, s183_10, s183_11, s183_12, s183_13, s183_14, s183_15, s183_16, s183_17, s183_18, s183_19, s183_20, s183_21, s183_22, s185, s187)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s185, const00000) = '1' then s188_0 <= s187; else s188_0 <= s183_0; end if;
     if equal(s185, const00001) = '1' then s188_1 <= s187; else s188_1 <= s183_1; end if;
     if equal(s185, const00010) = '1' then s188_2 <= s187; else s188_2 <= s183_2; end if;
     if equal(s185, const00011) = '1' then s188_3 <= s187; else s188_3 <= s183_3; end if;
     if equal(s185, const00100) = '1' then s188_4 <= s187; else s188_4 <= s183_4; end if;
     if equal(s185, const00101) = '1' then s188_5 <= s187; else s188_5 <= s183_5; end if;
     if equal(s185, const00110) = '1' then s188_6 <= s187; else s188_6 <= s183_6; end if;
     if equal(s185, const00111) = '1' then s188_7 <= s187; else s188_7 <= s183_7; end if;
     if equal(s185, const01000) = '1' then s188_8 <= s187; else s188_8 <= s183_8; end if;
     if equal(s185, const01001) = '1' then s188_9 <= s187; else s188_9 <= s183_9; end if;
     if equal(s185, const01010) = '1' then s188_10 <= s187; else s188_10 <= s183_10; end if;
     if equal(s185, const01011) = '1' then s188_11 <= s187; else s188_11 <= s183_11; end if;
     if equal(s185, const01100) = '1' then s188_12 <= s187; else s188_12 <= s183_12; end if;
     if equal(s185, const01101) = '1' then s188_13 <= s187; else s188_13 <= s183_13; end if;
     if equal(s185, const01110) = '1' then s188_14 <= s187; else s188_14 <= s183_14; end if;
     if equal(s185, const01111) = '1' then s188_15 <= s187; else s188_15 <= s183_15; end if;
     if equal(s185, const10000) = '1' then s188_16 <= s187; else s188_16 <= s183_16; end if;
     if equal(s185, const10001) = '1' then s188_17 <= s187; else s188_17 <= s183_17; end if;
     if equal(s185, const10010) = '1' then s188_18 <= s187; else s188_18 <= s183_18; end if;
     if equal(s185, const10011) = '1' then s188_19 <= s187; else s188_19 <= s183_19; end if;
     if equal(s185, const10100) = '1' then s188_20 <= s187; else s188_20 <= s183_20; end if;
     if equal(s185, const10101) = '1' then s188_21 <= s187; else s188_21 <= s183_21; end if;
     if equal(s185, const10110) = '1' then s188_22 <= s187; else s188_22 <= s183_22; end if;
   end process;

   s190 <= "01011";  -- constint module constint_11_157

   -- array reader array_reader_158
   process(s188_0, s188_1, s188_2, s188_3, s188_4, s188_5, s188_6, s188_7, s188_8, s188_9, s188_10, s188_11, s188_12, s188_13, s188_14, s188_15, s188_16, s188_17, s188_18, s188_19, s188_20, s188_21, s188_22, s190)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s190, const00000) = '1' ) then s191 <= s188_0; else
       if (equal(s190, const00001) = '1' ) then s191 <= s188_1; else
       if (equal(s190, const00010) = '1' ) then s191 <= s188_2; else
       if (equal(s190, const00011) = '1' ) then s191 <= s188_3; else
       if (equal(s190, const00100) = '1' ) then s191 <= s188_4; else
       if (equal(s190, const00101) = '1' ) then s191 <= s188_5; else
       if (equal(s190, const00110) = '1' ) then s191 <= s188_6; else
       if (equal(s190, const00111) = '1' ) then s191 <= s188_7; else
       if (equal(s190, const01000) = '1' ) then s191 <= s188_8; else
       if (equal(s190, const01001) = '1' ) then s191 <= s188_9; else
       if (equal(s190, const01010) = '1' ) then s191 <= s188_10; else
       if (equal(s190, const01011) = '1' ) then s191 <= s188_11; else
       if (equal(s190, const01100) = '1' ) then s191 <= s188_12; else
       if (equal(s190, const01101) = '1' ) then s191 <= s188_13; else
       if (equal(s190, const01110) = '1' ) then s191 <= s188_14; else
       if (equal(s190, const01111) = '1' ) then s191 <= s188_15; else
       if (equal(s190, const10000) = '1' ) then s191 <= s188_16; else
       if (equal(s190, const10001) = '1' ) then s191 <= s188_17; else
       if (equal(s190, const10010) = '1' ) then s191 <= s188_18; else
       if (equal(s190, const10011) = '1' ) then s191 <= s188_19; else
       if (equal(s190, const10100) = '1' ) then s191 <= s188_20; else
       if (equal(s190, const10101) = '1' ) then s191 <= s188_21; else
       s191 <= s188_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_159
   process(s133, s191, s189)
   begin
   if ( s133 = '1') then s192 <= s189; else s192 <= s191;
   end if;
   end process;

   -- array writer array_writer_160
   process(s188_0, s188_1, s188_2, s188_3, s188_4, s188_5, s188_6, s188_7, s188_8, s188_9, s188_10, s188_11, s188_12, s188_13, s188_14, s188_15, s188_16, s188_17, s188_18, s188_19, s188_20, s188_21, s188_22, s190, s192)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s190, const00000) = '1' then s193_0 <= s192; else s193_0 <= s188_0; end if;
     if equal(s190, const00001) = '1' then s193_1 <= s192; else s193_1 <= s188_1; end if;
     if equal(s190, const00010) = '1' then s193_2 <= s192; else s193_2 <= s188_2; end if;
     if equal(s190, const00011) = '1' then s193_3 <= s192; else s193_3 <= s188_3; end if;
     if equal(s190, const00100) = '1' then s193_4 <= s192; else s193_4 <= s188_4; end if;
     if equal(s190, const00101) = '1' then s193_5 <= s192; else s193_5 <= s188_5; end if;
     if equal(s190, const00110) = '1' then s193_6 <= s192; else s193_6 <= s188_6; end if;
     if equal(s190, const00111) = '1' then s193_7 <= s192; else s193_7 <= s188_7; end if;
     if equal(s190, const01000) = '1' then s193_8 <= s192; else s193_8 <= s188_8; end if;
     if equal(s190, const01001) = '1' then s193_9 <= s192; else s193_9 <= s188_9; end if;
     if equal(s190, const01010) = '1' then s193_10 <= s192; else s193_10 <= s188_10; end if;
     if equal(s190, const01011) = '1' then s193_11 <= s192; else s193_11 <= s188_11; end if;
     if equal(s190, const01100) = '1' then s193_12 <= s192; else s193_12 <= s188_12; end if;
     if equal(s190, const01101) = '1' then s193_13 <= s192; else s193_13 <= s188_13; end if;
     if equal(s190, const01110) = '1' then s193_14 <= s192; else s193_14 <= s188_14; end if;
     if equal(s190, const01111) = '1' then s193_15 <= s192; else s193_15 <= s188_15; end if;
     if equal(s190, const10000) = '1' then s193_16 <= s192; else s193_16 <= s188_16; end if;
     if equal(s190, const10001) = '1' then s193_17 <= s192; else s193_17 <= s188_17; end if;
     if equal(s190, const10010) = '1' then s193_18 <= s192; else s193_18 <= s188_18; end if;
     if equal(s190, const10011) = '1' then s193_19 <= s192; else s193_19 <= s188_19; end if;
     if equal(s190, const10100) = '1' then s193_20 <= s192; else s193_20 <= s188_20; end if;
     if equal(s190, const10101) = '1' then s193_21 <= s192; else s193_21 <= s188_21; end if;
     if equal(s190, const10110) = '1' then s193_22 <= s192; else s193_22 <= s188_22; end if;
   end process;

   s195 <= "01100";  -- constint module constint_12_161

   -- array reader array_reader_162
   process(s193_0, s193_1, s193_2, s193_3, s193_4, s193_5, s193_6, s193_7, s193_8, s193_9, s193_10, s193_11, s193_12, s193_13, s193_14, s193_15, s193_16, s193_17, s193_18, s193_19, s193_20, s193_21, s193_22, s195)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s195, const00000) = '1' ) then s196 <= s193_0; else
       if (equal(s195, const00001) = '1' ) then s196 <= s193_1; else
       if (equal(s195, const00010) = '1' ) then s196 <= s193_2; else
       if (equal(s195, const00011) = '1' ) then s196 <= s193_3; else
       if (equal(s195, const00100) = '1' ) then s196 <= s193_4; else
       if (equal(s195, const00101) = '1' ) then s196 <= s193_5; else
       if (equal(s195, const00110) = '1' ) then s196 <= s193_6; else
       if (equal(s195, const00111) = '1' ) then s196 <= s193_7; else
       if (equal(s195, const01000) = '1' ) then s196 <= s193_8; else
       if (equal(s195, const01001) = '1' ) then s196 <= s193_9; else
       if (equal(s195, const01010) = '1' ) then s196 <= s193_10; else
       if (equal(s195, const01011) = '1' ) then s196 <= s193_11; else
       if (equal(s195, const01100) = '1' ) then s196 <= s193_12; else
       if (equal(s195, const01101) = '1' ) then s196 <= s193_13; else
       if (equal(s195, const01110) = '1' ) then s196 <= s193_14; else
       if (equal(s195, const01111) = '1' ) then s196 <= s193_15; else
       if (equal(s195, const10000) = '1' ) then s196 <= s193_16; else
       if (equal(s195, const10001) = '1' ) then s196 <= s193_17; else
       if (equal(s195, const10010) = '1' ) then s196 <= s193_18; else
       if (equal(s195, const10011) = '1' ) then s196 <= s193_19; else
       if (equal(s195, const10100) = '1' ) then s196 <= s193_20; else
       if (equal(s195, const10101) = '1' ) then s196 <= s193_21; else
       s196 <= s193_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_163
   process(s133, s196, s194)
   begin
   if ( s133 = '1') then s197 <= s194; else s197 <= s196;
   end if;
   end process;

   -- array writer array_writer_164
   process(s193_0, s193_1, s193_2, s193_3, s193_4, s193_5, s193_6, s193_7, s193_8, s193_9, s193_10, s193_11, s193_12, s193_13, s193_14, s193_15, s193_16, s193_17, s193_18, s193_19, s193_20, s193_21, s193_22, s195, s197)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s195, const00000) = '1' then s198_0 <= s197; else s198_0 <= s193_0; end if;
     if equal(s195, const00001) = '1' then s198_1 <= s197; else s198_1 <= s193_1; end if;
     if equal(s195, const00010) = '1' then s198_2 <= s197; else s198_2 <= s193_2; end if;
     if equal(s195, const00011) = '1' then s198_3 <= s197; else s198_3 <= s193_3; end if;
     if equal(s195, const00100) = '1' then s198_4 <= s197; else s198_4 <= s193_4; end if;
     if equal(s195, const00101) = '1' then s198_5 <= s197; else s198_5 <= s193_5; end if;
     if equal(s195, const00110) = '1' then s198_6 <= s197; else s198_6 <= s193_6; end if;
     if equal(s195, const00111) = '1' then s198_7 <= s197; else s198_7 <= s193_7; end if;
     if equal(s195, const01000) = '1' then s198_8 <= s197; else s198_8 <= s193_8; end if;
     if equal(s195, const01001) = '1' then s198_9 <= s197; else s198_9 <= s193_9; end if;
     if equal(s195, const01010) = '1' then s198_10 <= s197; else s198_10 <= s193_10; end if;
     if equal(s195, const01011) = '1' then s198_11 <= s197; else s198_11 <= s193_11; end if;
     if equal(s195, const01100) = '1' then s198_12 <= s197; else s198_12 <= s193_12; end if;
     if equal(s195, const01101) = '1' then s198_13 <= s197; else s198_13 <= s193_13; end if;
     if equal(s195, const01110) = '1' then s198_14 <= s197; else s198_14 <= s193_14; end if;
     if equal(s195, const01111) = '1' then s198_15 <= s197; else s198_15 <= s193_15; end if;
     if equal(s195, const10000) = '1' then s198_16 <= s197; else s198_16 <= s193_16; end if;
     if equal(s195, const10001) = '1' then s198_17 <= s197; else s198_17 <= s193_17; end if;
     if equal(s195, const10010) = '1' then s198_18 <= s197; else s198_18 <= s193_18; end if;
     if equal(s195, const10011) = '1' then s198_19 <= s197; else s198_19 <= s193_19; end if;
     if equal(s195, const10100) = '1' then s198_20 <= s197; else s198_20 <= s193_20; end if;
     if equal(s195, const10101) = '1' then s198_21 <= s197; else s198_21 <= s193_21; end if;
     if equal(s195, const10110) = '1' then s198_22 <= s197; else s198_22 <= s193_22; end if;
   end process;

   s200 <= "01101";  -- constint module constint_13_165

   -- array reader array_reader_166
   process(s198_0, s198_1, s198_2, s198_3, s198_4, s198_5, s198_6, s198_7, s198_8, s198_9, s198_10, s198_11, s198_12, s198_13, s198_14, s198_15, s198_16, s198_17, s198_18, s198_19, s198_20, s198_21, s198_22, s200)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s200, const00000) = '1' ) then s201 <= s198_0; else
       if (equal(s200, const00001) = '1' ) then s201 <= s198_1; else
       if (equal(s200, const00010) = '1' ) then s201 <= s198_2; else
       if (equal(s200, const00011) = '1' ) then s201 <= s198_3; else
       if (equal(s200, const00100) = '1' ) then s201 <= s198_4; else
       if (equal(s200, const00101) = '1' ) then s201 <= s198_5; else
       if (equal(s200, const00110) = '1' ) then s201 <= s198_6; else
       if (equal(s200, const00111) = '1' ) then s201 <= s198_7; else
       if (equal(s200, const01000) = '1' ) then s201 <= s198_8; else
       if (equal(s200, const01001) = '1' ) then s201 <= s198_9; else
       if (equal(s200, const01010) = '1' ) then s201 <= s198_10; else
       if (equal(s200, const01011) = '1' ) then s201 <= s198_11; else
       if (equal(s200, const01100) = '1' ) then s201 <= s198_12; else
       if (equal(s200, const01101) = '1' ) then s201 <= s198_13; else
       if (equal(s200, const01110) = '1' ) then s201 <= s198_14; else
       if (equal(s200, const01111) = '1' ) then s201 <= s198_15; else
       if (equal(s200, const10000) = '1' ) then s201 <= s198_16; else
       if (equal(s200, const10001) = '1' ) then s201 <= s198_17; else
       if (equal(s200, const10010) = '1' ) then s201 <= s198_18; else
       if (equal(s200, const10011) = '1' ) then s201 <= s198_19; else
       if (equal(s200, const10100) = '1' ) then s201 <= s198_20; else
       if (equal(s200, const10101) = '1' ) then s201 <= s198_21; else
       s201 <= s198_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_167
   process(s133, s201, s199)
   begin
   if ( s133 = '1') then s202 <= s199; else s202 <= s201;
   end if;
   end process;

   -- array writer array_writer_168
   process(s198_0, s198_1, s198_2, s198_3, s198_4, s198_5, s198_6, s198_7, s198_8, s198_9, s198_10, s198_11, s198_12, s198_13, s198_14, s198_15, s198_16, s198_17, s198_18, s198_19, s198_20, s198_21, s198_22, s200, s202)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s200, const00000) = '1' then s203_0 <= s202; else s203_0 <= s198_0; end if;
     if equal(s200, const00001) = '1' then s203_1 <= s202; else s203_1 <= s198_1; end if;
     if equal(s200, const00010) = '1' then s203_2 <= s202; else s203_2 <= s198_2; end if;
     if equal(s200, const00011) = '1' then s203_3 <= s202; else s203_3 <= s198_3; end if;
     if equal(s200, const00100) = '1' then s203_4 <= s202; else s203_4 <= s198_4; end if;
     if equal(s200, const00101) = '1' then s203_5 <= s202; else s203_5 <= s198_5; end if;
     if equal(s200, const00110) = '1' then s203_6 <= s202; else s203_6 <= s198_6; end if;
     if equal(s200, const00111) = '1' then s203_7 <= s202; else s203_7 <= s198_7; end if;
     if equal(s200, const01000) = '1' then s203_8 <= s202; else s203_8 <= s198_8; end if;
     if equal(s200, const01001) = '1' then s203_9 <= s202; else s203_9 <= s198_9; end if;
     if equal(s200, const01010) = '1' then s203_10 <= s202; else s203_10 <= s198_10; end if;
     if equal(s200, const01011) = '1' then s203_11 <= s202; else s203_11 <= s198_11; end if;
     if equal(s200, const01100) = '1' then s203_12 <= s202; else s203_12 <= s198_12; end if;
     if equal(s200, const01101) = '1' then s203_13 <= s202; else s203_13 <= s198_13; end if;
     if equal(s200, const01110) = '1' then s203_14 <= s202; else s203_14 <= s198_14; end if;
     if equal(s200, const01111) = '1' then s203_15 <= s202; else s203_15 <= s198_15; end if;
     if equal(s200, const10000) = '1' then s203_16 <= s202; else s203_16 <= s198_16; end if;
     if equal(s200, const10001) = '1' then s203_17 <= s202; else s203_17 <= s198_17; end if;
     if equal(s200, const10010) = '1' then s203_18 <= s202; else s203_18 <= s198_18; end if;
     if equal(s200, const10011) = '1' then s203_19 <= s202; else s203_19 <= s198_19; end if;
     if equal(s200, const10100) = '1' then s203_20 <= s202; else s203_20 <= s198_20; end if;
     if equal(s200, const10101) = '1' then s203_21 <= s202; else s203_21 <= s198_21; end if;
     if equal(s200, const10110) = '1' then s203_22 <= s202; else s203_22 <= s198_22; end if;
   end process;

   s205 <= "01110";  -- constint module constint_14_169

   -- array reader array_reader_170
   process(s203_0, s203_1, s203_2, s203_3, s203_4, s203_5, s203_6, s203_7, s203_8, s203_9, s203_10, s203_11, s203_12, s203_13, s203_14, s203_15, s203_16, s203_17, s203_18, s203_19, s203_20, s203_21, s203_22, s205)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s205, const00000) = '1' ) then s206 <= s203_0; else
       if (equal(s205, const00001) = '1' ) then s206 <= s203_1; else
       if (equal(s205, const00010) = '1' ) then s206 <= s203_2; else
       if (equal(s205, const00011) = '1' ) then s206 <= s203_3; else
       if (equal(s205, const00100) = '1' ) then s206 <= s203_4; else
       if (equal(s205, const00101) = '1' ) then s206 <= s203_5; else
       if (equal(s205, const00110) = '1' ) then s206 <= s203_6; else
       if (equal(s205, const00111) = '1' ) then s206 <= s203_7; else
       if (equal(s205, const01000) = '1' ) then s206 <= s203_8; else
       if (equal(s205, const01001) = '1' ) then s206 <= s203_9; else
       if (equal(s205, const01010) = '1' ) then s206 <= s203_10; else
       if (equal(s205, const01011) = '1' ) then s206 <= s203_11; else
       if (equal(s205, const01100) = '1' ) then s206 <= s203_12; else
       if (equal(s205, const01101) = '1' ) then s206 <= s203_13; else
       if (equal(s205, const01110) = '1' ) then s206 <= s203_14; else
       if (equal(s205, const01111) = '1' ) then s206 <= s203_15; else
       if (equal(s205, const10000) = '1' ) then s206 <= s203_16; else
       if (equal(s205, const10001) = '1' ) then s206 <= s203_17; else
       if (equal(s205, const10010) = '1' ) then s206 <= s203_18; else
       if (equal(s205, const10011) = '1' ) then s206 <= s203_19; else
       if (equal(s205, const10100) = '1' ) then s206 <= s203_20; else
       if (equal(s205, const10101) = '1' ) then s206 <= s203_21; else
       s206 <= s203_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_171
   process(s133, s206, s204)
   begin
   if ( s133 = '1') then s207 <= s204; else s207 <= s206;
   end if;
   end process;

   -- array writer array_writer_172
   process(s203_0, s203_1, s203_2, s203_3, s203_4, s203_5, s203_6, s203_7, s203_8, s203_9, s203_10, s203_11, s203_12, s203_13, s203_14, s203_15, s203_16, s203_17, s203_18, s203_19, s203_20, s203_21, s203_22, s205, s207)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s205, const00000) = '1' then s208_0 <= s207; else s208_0 <= s203_0; end if;
     if equal(s205, const00001) = '1' then s208_1 <= s207; else s208_1 <= s203_1; end if;
     if equal(s205, const00010) = '1' then s208_2 <= s207; else s208_2 <= s203_2; end if;
     if equal(s205, const00011) = '1' then s208_3 <= s207; else s208_3 <= s203_3; end if;
     if equal(s205, const00100) = '1' then s208_4 <= s207; else s208_4 <= s203_4; end if;
     if equal(s205, const00101) = '1' then s208_5 <= s207; else s208_5 <= s203_5; end if;
     if equal(s205, const00110) = '1' then s208_6 <= s207; else s208_6 <= s203_6; end if;
     if equal(s205, const00111) = '1' then s208_7 <= s207; else s208_7 <= s203_7; end if;
     if equal(s205, const01000) = '1' then s208_8 <= s207; else s208_8 <= s203_8; end if;
     if equal(s205, const01001) = '1' then s208_9 <= s207; else s208_9 <= s203_9; end if;
     if equal(s205, const01010) = '1' then s208_10 <= s207; else s208_10 <= s203_10; end if;
     if equal(s205, const01011) = '1' then s208_11 <= s207; else s208_11 <= s203_11; end if;
     if equal(s205, const01100) = '1' then s208_12 <= s207; else s208_12 <= s203_12; end if;
     if equal(s205, const01101) = '1' then s208_13 <= s207; else s208_13 <= s203_13; end if;
     if equal(s205, const01110) = '1' then s208_14 <= s207; else s208_14 <= s203_14; end if;
     if equal(s205, const01111) = '1' then s208_15 <= s207; else s208_15 <= s203_15; end if;
     if equal(s205, const10000) = '1' then s208_16 <= s207; else s208_16 <= s203_16; end if;
     if equal(s205, const10001) = '1' then s208_17 <= s207; else s208_17 <= s203_17; end if;
     if equal(s205, const10010) = '1' then s208_18 <= s207; else s208_18 <= s203_18; end if;
     if equal(s205, const10011) = '1' then s208_19 <= s207; else s208_19 <= s203_19; end if;
     if equal(s205, const10100) = '1' then s208_20 <= s207; else s208_20 <= s203_20; end if;
     if equal(s205, const10101) = '1' then s208_21 <= s207; else s208_21 <= s203_21; end if;
     if equal(s205, const10110) = '1' then s208_22 <= s207; else s208_22 <= s203_22; end if;
   end process;

   s210 <= "01111";  -- constint module constint_15_173

   -- array reader array_reader_174
   process(s208_0, s208_1, s208_2, s208_3, s208_4, s208_5, s208_6, s208_7, s208_8, s208_9, s208_10, s208_11, s208_12, s208_13, s208_14, s208_15, s208_16, s208_17, s208_18, s208_19, s208_20, s208_21, s208_22, s210)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s210, const00000) = '1' ) then s211 <= s208_0; else
       if (equal(s210, const00001) = '1' ) then s211 <= s208_1; else
       if (equal(s210, const00010) = '1' ) then s211 <= s208_2; else
       if (equal(s210, const00011) = '1' ) then s211 <= s208_3; else
       if (equal(s210, const00100) = '1' ) then s211 <= s208_4; else
       if (equal(s210, const00101) = '1' ) then s211 <= s208_5; else
       if (equal(s210, const00110) = '1' ) then s211 <= s208_6; else
       if (equal(s210, const00111) = '1' ) then s211 <= s208_7; else
       if (equal(s210, const01000) = '1' ) then s211 <= s208_8; else
       if (equal(s210, const01001) = '1' ) then s211 <= s208_9; else
       if (equal(s210, const01010) = '1' ) then s211 <= s208_10; else
       if (equal(s210, const01011) = '1' ) then s211 <= s208_11; else
       if (equal(s210, const01100) = '1' ) then s211 <= s208_12; else
       if (equal(s210, const01101) = '1' ) then s211 <= s208_13; else
       if (equal(s210, const01110) = '1' ) then s211 <= s208_14; else
       if (equal(s210, const01111) = '1' ) then s211 <= s208_15; else
       if (equal(s210, const10000) = '1' ) then s211 <= s208_16; else
       if (equal(s210, const10001) = '1' ) then s211 <= s208_17; else
       if (equal(s210, const10010) = '1' ) then s211 <= s208_18; else
       if (equal(s210, const10011) = '1' ) then s211 <= s208_19; else
       if (equal(s210, const10100) = '1' ) then s211 <= s208_20; else
       if (equal(s210, const10101) = '1' ) then s211 <= s208_21; else
       s211 <= s208_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_175
   process(s133, s211, s209)
   begin
   if ( s133 = '1') then s212 <= s209; else s212 <= s211;
   end if;
   end process;

   -- array writer array_writer_176
   process(s208_0, s208_1, s208_2, s208_3, s208_4, s208_5, s208_6, s208_7, s208_8, s208_9, s208_10, s208_11, s208_12, s208_13, s208_14, s208_15, s208_16, s208_17, s208_18, s208_19, s208_20, s208_21, s208_22, s210, s212)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s210, const00000) = '1' then s213_0 <= s212; else s213_0 <= s208_0; end if;
     if equal(s210, const00001) = '1' then s213_1 <= s212; else s213_1 <= s208_1; end if;
     if equal(s210, const00010) = '1' then s213_2 <= s212; else s213_2 <= s208_2; end if;
     if equal(s210, const00011) = '1' then s213_3 <= s212; else s213_3 <= s208_3; end if;
     if equal(s210, const00100) = '1' then s213_4 <= s212; else s213_4 <= s208_4; end if;
     if equal(s210, const00101) = '1' then s213_5 <= s212; else s213_5 <= s208_5; end if;
     if equal(s210, const00110) = '1' then s213_6 <= s212; else s213_6 <= s208_6; end if;
     if equal(s210, const00111) = '1' then s213_7 <= s212; else s213_7 <= s208_7; end if;
     if equal(s210, const01000) = '1' then s213_8 <= s212; else s213_8 <= s208_8; end if;
     if equal(s210, const01001) = '1' then s213_9 <= s212; else s213_9 <= s208_9; end if;
     if equal(s210, const01010) = '1' then s213_10 <= s212; else s213_10 <= s208_10; end if;
     if equal(s210, const01011) = '1' then s213_11 <= s212; else s213_11 <= s208_11; end if;
     if equal(s210, const01100) = '1' then s213_12 <= s212; else s213_12 <= s208_12; end if;
     if equal(s210, const01101) = '1' then s213_13 <= s212; else s213_13 <= s208_13; end if;
     if equal(s210, const01110) = '1' then s213_14 <= s212; else s213_14 <= s208_14; end if;
     if equal(s210, const01111) = '1' then s213_15 <= s212; else s213_15 <= s208_15; end if;
     if equal(s210, const10000) = '1' then s213_16 <= s212; else s213_16 <= s208_16; end if;
     if equal(s210, const10001) = '1' then s213_17 <= s212; else s213_17 <= s208_17; end if;
     if equal(s210, const10010) = '1' then s213_18 <= s212; else s213_18 <= s208_18; end if;
     if equal(s210, const10011) = '1' then s213_19 <= s212; else s213_19 <= s208_19; end if;
     if equal(s210, const10100) = '1' then s213_20 <= s212; else s213_20 <= s208_20; end if;
     if equal(s210, const10101) = '1' then s213_21 <= s212; else s213_21 <= s208_21; end if;
     if equal(s210, const10110) = '1' then s213_22 <= s212; else s213_22 <= s208_22; end if;
   end process;

   s215 <= "10000";  -- constint module constint_16_177

   -- array reader array_reader_178
   process(s213_0, s213_1, s213_2, s213_3, s213_4, s213_5, s213_6, s213_7, s213_8, s213_9, s213_10, s213_11, s213_12, s213_13, s213_14, s213_15, s213_16, s213_17, s213_18, s213_19, s213_20, s213_21, s213_22, s215)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s215, const00000) = '1' ) then s216 <= s213_0; else
       if (equal(s215, const00001) = '1' ) then s216 <= s213_1; else
       if (equal(s215, const00010) = '1' ) then s216 <= s213_2; else
       if (equal(s215, const00011) = '1' ) then s216 <= s213_3; else
       if (equal(s215, const00100) = '1' ) then s216 <= s213_4; else
       if (equal(s215, const00101) = '1' ) then s216 <= s213_5; else
       if (equal(s215, const00110) = '1' ) then s216 <= s213_6; else
       if (equal(s215, const00111) = '1' ) then s216 <= s213_7; else
       if (equal(s215, const01000) = '1' ) then s216 <= s213_8; else
       if (equal(s215, const01001) = '1' ) then s216 <= s213_9; else
       if (equal(s215, const01010) = '1' ) then s216 <= s213_10; else
       if (equal(s215, const01011) = '1' ) then s216 <= s213_11; else
       if (equal(s215, const01100) = '1' ) then s216 <= s213_12; else
       if (equal(s215, const01101) = '1' ) then s216 <= s213_13; else
       if (equal(s215, const01110) = '1' ) then s216 <= s213_14; else
       if (equal(s215, const01111) = '1' ) then s216 <= s213_15; else
       if (equal(s215, const10000) = '1' ) then s216 <= s213_16; else
       if (equal(s215, const10001) = '1' ) then s216 <= s213_17; else
       if (equal(s215, const10010) = '1' ) then s216 <= s213_18; else
       if (equal(s215, const10011) = '1' ) then s216 <= s213_19; else
       if (equal(s215, const10100) = '1' ) then s216 <= s213_20; else
       if (equal(s215, const10101) = '1' ) then s216 <= s213_21; else
       s216 <= s213_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_179
   process(s133, s216, s214)
   begin
   if ( s133 = '1') then s217 <= s214; else s217 <= s216;
   end if;
   end process;

   -- array writer array_writer_180
   process(s213_0, s213_1, s213_2, s213_3, s213_4, s213_5, s213_6, s213_7, s213_8, s213_9, s213_10, s213_11, s213_12, s213_13, s213_14, s213_15, s213_16, s213_17, s213_18, s213_19, s213_20, s213_21, s213_22, s215, s217)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s215, const00000) = '1' then s218_0 <= s217; else s218_0 <= s213_0; end if;
     if equal(s215, const00001) = '1' then s218_1 <= s217; else s218_1 <= s213_1; end if;
     if equal(s215, const00010) = '1' then s218_2 <= s217; else s218_2 <= s213_2; end if;
     if equal(s215, const00011) = '1' then s218_3 <= s217; else s218_3 <= s213_3; end if;
     if equal(s215, const00100) = '1' then s218_4 <= s217; else s218_4 <= s213_4; end if;
     if equal(s215, const00101) = '1' then s218_5 <= s217; else s218_5 <= s213_5; end if;
     if equal(s215, const00110) = '1' then s218_6 <= s217; else s218_6 <= s213_6; end if;
     if equal(s215, const00111) = '1' then s218_7 <= s217; else s218_7 <= s213_7; end if;
     if equal(s215, const01000) = '1' then s218_8 <= s217; else s218_8 <= s213_8; end if;
     if equal(s215, const01001) = '1' then s218_9 <= s217; else s218_9 <= s213_9; end if;
     if equal(s215, const01010) = '1' then s218_10 <= s217; else s218_10 <= s213_10; end if;
     if equal(s215, const01011) = '1' then s218_11 <= s217; else s218_11 <= s213_11; end if;
     if equal(s215, const01100) = '1' then s218_12 <= s217; else s218_12 <= s213_12; end if;
     if equal(s215, const01101) = '1' then s218_13 <= s217; else s218_13 <= s213_13; end if;
     if equal(s215, const01110) = '1' then s218_14 <= s217; else s218_14 <= s213_14; end if;
     if equal(s215, const01111) = '1' then s218_15 <= s217; else s218_15 <= s213_15; end if;
     if equal(s215, const10000) = '1' then s218_16 <= s217; else s218_16 <= s213_16; end if;
     if equal(s215, const10001) = '1' then s218_17 <= s217; else s218_17 <= s213_17; end if;
     if equal(s215, const10010) = '1' then s218_18 <= s217; else s218_18 <= s213_18; end if;
     if equal(s215, const10011) = '1' then s218_19 <= s217; else s218_19 <= s213_19; end if;
     if equal(s215, const10100) = '1' then s218_20 <= s217; else s218_20 <= s213_20; end if;
     if equal(s215, const10101) = '1' then s218_21 <= s217; else s218_21 <= s213_21; end if;
     if equal(s215, const10110) = '1' then s218_22 <= s217; else s218_22 <= s213_22; end if;
   end process;

   s220 <= "10001";  -- constint module constint_17_181

   -- array reader array_reader_182
   process(s218_0, s218_1, s218_2, s218_3, s218_4, s218_5, s218_6, s218_7, s218_8, s218_9, s218_10, s218_11, s218_12, s218_13, s218_14, s218_15, s218_16, s218_17, s218_18, s218_19, s218_20, s218_21, s218_22, s220)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s220, const00000) = '1' ) then s221 <= s218_0; else
       if (equal(s220, const00001) = '1' ) then s221 <= s218_1; else
       if (equal(s220, const00010) = '1' ) then s221 <= s218_2; else
       if (equal(s220, const00011) = '1' ) then s221 <= s218_3; else
       if (equal(s220, const00100) = '1' ) then s221 <= s218_4; else
       if (equal(s220, const00101) = '1' ) then s221 <= s218_5; else
       if (equal(s220, const00110) = '1' ) then s221 <= s218_6; else
       if (equal(s220, const00111) = '1' ) then s221 <= s218_7; else
       if (equal(s220, const01000) = '1' ) then s221 <= s218_8; else
       if (equal(s220, const01001) = '1' ) then s221 <= s218_9; else
       if (equal(s220, const01010) = '1' ) then s221 <= s218_10; else
       if (equal(s220, const01011) = '1' ) then s221 <= s218_11; else
       if (equal(s220, const01100) = '1' ) then s221 <= s218_12; else
       if (equal(s220, const01101) = '1' ) then s221 <= s218_13; else
       if (equal(s220, const01110) = '1' ) then s221 <= s218_14; else
       if (equal(s220, const01111) = '1' ) then s221 <= s218_15; else
       if (equal(s220, const10000) = '1' ) then s221 <= s218_16; else
       if (equal(s220, const10001) = '1' ) then s221 <= s218_17; else
       if (equal(s220, const10010) = '1' ) then s221 <= s218_18; else
       if (equal(s220, const10011) = '1' ) then s221 <= s218_19; else
       if (equal(s220, const10100) = '1' ) then s221 <= s218_20; else
       if (equal(s220, const10101) = '1' ) then s221 <= s218_21; else
       s221 <= s218_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_183
   process(s133, s221, s219)
   begin
   if ( s133 = '1') then s222 <= s219; else s222 <= s221;
   end if;
   end process;

   -- array writer array_writer_184
   process(s218_0, s218_1, s218_2, s218_3, s218_4, s218_5, s218_6, s218_7, s218_8, s218_9, s218_10, s218_11, s218_12, s218_13, s218_14, s218_15, s218_16, s218_17, s218_18, s218_19, s218_20, s218_21, s218_22, s220, s222)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s220, const00000) = '1' then s223_0 <= s222; else s223_0 <= s218_0; end if;
     if equal(s220, const00001) = '1' then s223_1 <= s222; else s223_1 <= s218_1; end if;
     if equal(s220, const00010) = '1' then s223_2 <= s222; else s223_2 <= s218_2; end if;
     if equal(s220, const00011) = '1' then s223_3 <= s222; else s223_3 <= s218_3; end if;
     if equal(s220, const00100) = '1' then s223_4 <= s222; else s223_4 <= s218_4; end if;
     if equal(s220, const00101) = '1' then s223_5 <= s222; else s223_5 <= s218_5; end if;
     if equal(s220, const00110) = '1' then s223_6 <= s222; else s223_6 <= s218_6; end if;
     if equal(s220, const00111) = '1' then s223_7 <= s222; else s223_7 <= s218_7; end if;
     if equal(s220, const01000) = '1' then s223_8 <= s222; else s223_8 <= s218_8; end if;
     if equal(s220, const01001) = '1' then s223_9 <= s222; else s223_9 <= s218_9; end if;
     if equal(s220, const01010) = '1' then s223_10 <= s222; else s223_10 <= s218_10; end if;
     if equal(s220, const01011) = '1' then s223_11 <= s222; else s223_11 <= s218_11; end if;
     if equal(s220, const01100) = '1' then s223_12 <= s222; else s223_12 <= s218_12; end if;
     if equal(s220, const01101) = '1' then s223_13 <= s222; else s223_13 <= s218_13; end if;
     if equal(s220, const01110) = '1' then s223_14 <= s222; else s223_14 <= s218_14; end if;
     if equal(s220, const01111) = '1' then s223_15 <= s222; else s223_15 <= s218_15; end if;
     if equal(s220, const10000) = '1' then s223_16 <= s222; else s223_16 <= s218_16; end if;
     if equal(s220, const10001) = '1' then s223_17 <= s222; else s223_17 <= s218_17; end if;
     if equal(s220, const10010) = '1' then s223_18 <= s222; else s223_18 <= s218_18; end if;
     if equal(s220, const10011) = '1' then s223_19 <= s222; else s223_19 <= s218_19; end if;
     if equal(s220, const10100) = '1' then s223_20 <= s222; else s223_20 <= s218_20; end if;
     if equal(s220, const10101) = '1' then s223_21 <= s222; else s223_21 <= s218_21; end if;
     if equal(s220, const10110) = '1' then s223_22 <= s222; else s223_22 <= s218_22; end if;
   end process;

   s225 <= "10010";  -- constint module constint_18_185

   -- array reader array_reader_186
   process(s223_0, s223_1, s223_2, s223_3, s223_4, s223_5, s223_6, s223_7, s223_8, s223_9, s223_10, s223_11, s223_12, s223_13, s223_14, s223_15, s223_16, s223_17, s223_18, s223_19, s223_20, s223_21, s223_22, s225)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s225, const00000) = '1' ) then s226 <= s223_0; else
       if (equal(s225, const00001) = '1' ) then s226 <= s223_1; else
       if (equal(s225, const00010) = '1' ) then s226 <= s223_2; else
       if (equal(s225, const00011) = '1' ) then s226 <= s223_3; else
       if (equal(s225, const00100) = '1' ) then s226 <= s223_4; else
       if (equal(s225, const00101) = '1' ) then s226 <= s223_5; else
       if (equal(s225, const00110) = '1' ) then s226 <= s223_6; else
       if (equal(s225, const00111) = '1' ) then s226 <= s223_7; else
       if (equal(s225, const01000) = '1' ) then s226 <= s223_8; else
       if (equal(s225, const01001) = '1' ) then s226 <= s223_9; else
       if (equal(s225, const01010) = '1' ) then s226 <= s223_10; else
       if (equal(s225, const01011) = '1' ) then s226 <= s223_11; else
       if (equal(s225, const01100) = '1' ) then s226 <= s223_12; else
       if (equal(s225, const01101) = '1' ) then s226 <= s223_13; else
       if (equal(s225, const01110) = '1' ) then s226 <= s223_14; else
       if (equal(s225, const01111) = '1' ) then s226 <= s223_15; else
       if (equal(s225, const10000) = '1' ) then s226 <= s223_16; else
       if (equal(s225, const10001) = '1' ) then s226 <= s223_17; else
       if (equal(s225, const10010) = '1' ) then s226 <= s223_18; else
       if (equal(s225, const10011) = '1' ) then s226 <= s223_19; else
       if (equal(s225, const10100) = '1' ) then s226 <= s223_20; else
       if (equal(s225, const10101) = '1' ) then s226 <= s223_21; else
       s226 <= s223_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_187
   process(s133, s226, s224)
   begin
   if ( s133 = '1') then s227 <= s224; else s227 <= s226;
   end if;
   end process;

   -- array writer array_writer_188
   process(s223_0, s223_1, s223_2, s223_3, s223_4, s223_5, s223_6, s223_7, s223_8, s223_9, s223_10, s223_11, s223_12, s223_13, s223_14, s223_15, s223_16, s223_17, s223_18, s223_19, s223_20, s223_21, s223_22, s225, s227)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s225, const00000) = '1' then s228_0 <= s227; else s228_0 <= s223_0; end if;
     if equal(s225, const00001) = '1' then s228_1 <= s227; else s228_1 <= s223_1; end if;
     if equal(s225, const00010) = '1' then s228_2 <= s227; else s228_2 <= s223_2; end if;
     if equal(s225, const00011) = '1' then s228_3 <= s227; else s228_3 <= s223_3; end if;
     if equal(s225, const00100) = '1' then s228_4 <= s227; else s228_4 <= s223_4; end if;
     if equal(s225, const00101) = '1' then s228_5 <= s227; else s228_5 <= s223_5; end if;
     if equal(s225, const00110) = '1' then s228_6 <= s227; else s228_6 <= s223_6; end if;
     if equal(s225, const00111) = '1' then s228_7 <= s227; else s228_7 <= s223_7; end if;
     if equal(s225, const01000) = '1' then s228_8 <= s227; else s228_8 <= s223_8; end if;
     if equal(s225, const01001) = '1' then s228_9 <= s227; else s228_9 <= s223_9; end if;
     if equal(s225, const01010) = '1' then s228_10 <= s227; else s228_10 <= s223_10; end if;
     if equal(s225, const01011) = '1' then s228_11 <= s227; else s228_11 <= s223_11; end if;
     if equal(s225, const01100) = '1' then s228_12 <= s227; else s228_12 <= s223_12; end if;
     if equal(s225, const01101) = '1' then s228_13 <= s227; else s228_13 <= s223_13; end if;
     if equal(s225, const01110) = '1' then s228_14 <= s227; else s228_14 <= s223_14; end if;
     if equal(s225, const01111) = '1' then s228_15 <= s227; else s228_15 <= s223_15; end if;
     if equal(s225, const10000) = '1' then s228_16 <= s227; else s228_16 <= s223_16; end if;
     if equal(s225, const10001) = '1' then s228_17 <= s227; else s228_17 <= s223_17; end if;
     if equal(s225, const10010) = '1' then s228_18 <= s227; else s228_18 <= s223_18; end if;
     if equal(s225, const10011) = '1' then s228_19 <= s227; else s228_19 <= s223_19; end if;
     if equal(s225, const10100) = '1' then s228_20 <= s227; else s228_20 <= s223_20; end if;
     if equal(s225, const10101) = '1' then s228_21 <= s227; else s228_21 <= s223_21; end if;
     if equal(s225, const10110) = '1' then s228_22 <= s227; else s228_22 <= s223_22; end if;
   end process;

   s230 <= "10011";  -- constint module constint_19_189

   -- array reader array_reader_190
   process(s228_0, s228_1, s228_2, s228_3, s228_4, s228_5, s228_6, s228_7, s228_8, s228_9, s228_10, s228_11, s228_12, s228_13, s228_14, s228_15, s228_16, s228_17, s228_18, s228_19, s228_20, s228_21, s228_22, s230)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s230, const00000) = '1' ) then s231 <= s228_0; else
       if (equal(s230, const00001) = '1' ) then s231 <= s228_1; else
       if (equal(s230, const00010) = '1' ) then s231 <= s228_2; else
       if (equal(s230, const00011) = '1' ) then s231 <= s228_3; else
       if (equal(s230, const00100) = '1' ) then s231 <= s228_4; else
       if (equal(s230, const00101) = '1' ) then s231 <= s228_5; else
       if (equal(s230, const00110) = '1' ) then s231 <= s228_6; else
       if (equal(s230, const00111) = '1' ) then s231 <= s228_7; else
       if (equal(s230, const01000) = '1' ) then s231 <= s228_8; else
       if (equal(s230, const01001) = '1' ) then s231 <= s228_9; else
       if (equal(s230, const01010) = '1' ) then s231 <= s228_10; else
       if (equal(s230, const01011) = '1' ) then s231 <= s228_11; else
       if (equal(s230, const01100) = '1' ) then s231 <= s228_12; else
       if (equal(s230, const01101) = '1' ) then s231 <= s228_13; else
       if (equal(s230, const01110) = '1' ) then s231 <= s228_14; else
       if (equal(s230, const01111) = '1' ) then s231 <= s228_15; else
       if (equal(s230, const10000) = '1' ) then s231 <= s228_16; else
       if (equal(s230, const10001) = '1' ) then s231 <= s228_17; else
       if (equal(s230, const10010) = '1' ) then s231 <= s228_18; else
       if (equal(s230, const10011) = '1' ) then s231 <= s228_19; else
       if (equal(s230, const10100) = '1' ) then s231 <= s228_20; else
       if (equal(s230, const10101) = '1' ) then s231 <= s228_21; else
       s231 <= s228_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_191
   process(s133, s231, s229)
   begin
   if ( s133 = '1') then s232 <= s229; else s232 <= s231;
   end if;
   end process;

   -- array writer array_writer_192
   process(s228_0, s228_1, s228_2, s228_3, s228_4, s228_5, s228_6, s228_7, s228_8, s228_9, s228_10, s228_11, s228_12, s228_13, s228_14, s228_15, s228_16, s228_17, s228_18, s228_19, s228_20, s228_21, s228_22, s230, s232)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s230, const00000) = '1' then s233_0 <= s232; else s233_0 <= s228_0; end if;
     if equal(s230, const00001) = '1' then s233_1 <= s232; else s233_1 <= s228_1; end if;
     if equal(s230, const00010) = '1' then s233_2 <= s232; else s233_2 <= s228_2; end if;
     if equal(s230, const00011) = '1' then s233_3 <= s232; else s233_3 <= s228_3; end if;
     if equal(s230, const00100) = '1' then s233_4 <= s232; else s233_4 <= s228_4; end if;
     if equal(s230, const00101) = '1' then s233_5 <= s232; else s233_5 <= s228_5; end if;
     if equal(s230, const00110) = '1' then s233_6 <= s232; else s233_6 <= s228_6; end if;
     if equal(s230, const00111) = '1' then s233_7 <= s232; else s233_7 <= s228_7; end if;
     if equal(s230, const01000) = '1' then s233_8 <= s232; else s233_8 <= s228_8; end if;
     if equal(s230, const01001) = '1' then s233_9 <= s232; else s233_9 <= s228_9; end if;
     if equal(s230, const01010) = '1' then s233_10 <= s232; else s233_10 <= s228_10; end if;
     if equal(s230, const01011) = '1' then s233_11 <= s232; else s233_11 <= s228_11; end if;
     if equal(s230, const01100) = '1' then s233_12 <= s232; else s233_12 <= s228_12; end if;
     if equal(s230, const01101) = '1' then s233_13 <= s232; else s233_13 <= s228_13; end if;
     if equal(s230, const01110) = '1' then s233_14 <= s232; else s233_14 <= s228_14; end if;
     if equal(s230, const01111) = '1' then s233_15 <= s232; else s233_15 <= s228_15; end if;
     if equal(s230, const10000) = '1' then s233_16 <= s232; else s233_16 <= s228_16; end if;
     if equal(s230, const10001) = '1' then s233_17 <= s232; else s233_17 <= s228_17; end if;
     if equal(s230, const10010) = '1' then s233_18 <= s232; else s233_18 <= s228_18; end if;
     if equal(s230, const10011) = '1' then s233_19 <= s232; else s233_19 <= s228_19; end if;
     if equal(s230, const10100) = '1' then s233_20 <= s232; else s233_20 <= s228_20; end if;
     if equal(s230, const10101) = '1' then s233_21 <= s232; else s233_21 <= s228_21; end if;
     if equal(s230, const10110) = '1' then s233_22 <= s232; else s233_22 <= s228_22; end if;
   end process;

   s235 <= "10100";  -- constint module constint_20_193

   -- array reader array_reader_194
   process(s233_0, s233_1, s233_2, s233_3, s233_4, s233_5, s233_6, s233_7, s233_8, s233_9, s233_10, s233_11, s233_12, s233_13, s233_14, s233_15, s233_16, s233_17, s233_18, s233_19, s233_20, s233_21, s233_22, s235)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s235, const00000) = '1' ) then s236 <= s233_0; else
       if (equal(s235, const00001) = '1' ) then s236 <= s233_1; else
       if (equal(s235, const00010) = '1' ) then s236 <= s233_2; else
       if (equal(s235, const00011) = '1' ) then s236 <= s233_3; else
       if (equal(s235, const00100) = '1' ) then s236 <= s233_4; else
       if (equal(s235, const00101) = '1' ) then s236 <= s233_5; else
       if (equal(s235, const00110) = '1' ) then s236 <= s233_6; else
       if (equal(s235, const00111) = '1' ) then s236 <= s233_7; else
       if (equal(s235, const01000) = '1' ) then s236 <= s233_8; else
       if (equal(s235, const01001) = '1' ) then s236 <= s233_9; else
       if (equal(s235, const01010) = '1' ) then s236 <= s233_10; else
       if (equal(s235, const01011) = '1' ) then s236 <= s233_11; else
       if (equal(s235, const01100) = '1' ) then s236 <= s233_12; else
       if (equal(s235, const01101) = '1' ) then s236 <= s233_13; else
       if (equal(s235, const01110) = '1' ) then s236 <= s233_14; else
       if (equal(s235, const01111) = '1' ) then s236 <= s233_15; else
       if (equal(s235, const10000) = '1' ) then s236 <= s233_16; else
       if (equal(s235, const10001) = '1' ) then s236 <= s233_17; else
       if (equal(s235, const10010) = '1' ) then s236 <= s233_18; else
       if (equal(s235, const10011) = '1' ) then s236 <= s233_19; else
       if (equal(s235, const10100) = '1' ) then s236 <= s233_20; else
       if (equal(s235, const10101) = '1' ) then s236 <= s233_21; else
       s236 <= s233_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_195
   process(s133, s236, s234)
   begin
   if ( s133 = '1') then s237 <= s234; else s237 <= s236;
   end if;
   end process;

   -- array writer array_writer_196
   process(s233_0, s233_1, s233_2, s233_3, s233_4, s233_5, s233_6, s233_7, s233_8, s233_9, s233_10, s233_11, s233_12, s233_13, s233_14, s233_15, s233_16, s233_17, s233_18, s233_19, s233_20, s233_21, s233_22, s235, s237)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s235, const00000) = '1' then s238_0 <= s237; else s238_0 <= s233_0; end if;
     if equal(s235, const00001) = '1' then s238_1 <= s237; else s238_1 <= s233_1; end if;
     if equal(s235, const00010) = '1' then s238_2 <= s237; else s238_2 <= s233_2; end if;
     if equal(s235, const00011) = '1' then s238_3 <= s237; else s238_3 <= s233_3; end if;
     if equal(s235, const00100) = '1' then s238_4 <= s237; else s238_4 <= s233_4; end if;
     if equal(s235, const00101) = '1' then s238_5 <= s237; else s238_5 <= s233_5; end if;
     if equal(s235, const00110) = '1' then s238_6 <= s237; else s238_6 <= s233_6; end if;
     if equal(s235, const00111) = '1' then s238_7 <= s237; else s238_7 <= s233_7; end if;
     if equal(s235, const01000) = '1' then s238_8 <= s237; else s238_8 <= s233_8; end if;
     if equal(s235, const01001) = '1' then s238_9 <= s237; else s238_9 <= s233_9; end if;
     if equal(s235, const01010) = '1' then s238_10 <= s237; else s238_10 <= s233_10; end if;
     if equal(s235, const01011) = '1' then s238_11 <= s237; else s238_11 <= s233_11; end if;
     if equal(s235, const01100) = '1' then s238_12 <= s237; else s238_12 <= s233_12; end if;
     if equal(s235, const01101) = '1' then s238_13 <= s237; else s238_13 <= s233_13; end if;
     if equal(s235, const01110) = '1' then s238_14 <= s237; else s238_14 <= s233_14; end if;
     if equal(s235, const01111) = '1' then s238_15 <= s237; else s238_15 <= s233_15; end if;
     if equal(s235, const10000) = '1' then s238_16 <= s237; else s238_16 <= s233_16; end if;
     if equal(s235, const10001) = '1' then s238_17 <= s237; else s238_17 <= s233_17; end if;
     if equal(s235, const10010) = '1' then s238_18 <= s237; else s238_18 <= s233_18; end if;
     if equal(s235, const10011) = '1' then s238_19 <= s237; else s238_19 <= s233_19; end if;
     if equal(s235, const10100) = '1' then s238_20 <= s237; else s238_20 <= s233_20; end if;
     if equal(s235, const10101) = '1' then s238_21 <= s237; else s238_21 <= s233_21; end if;
     if equal(s235, const10110) = '1' then s238_22 <= s237; else s238_22 <= s233_22; end if;
   end process;

   s240 <= "10101";  -- constint module constint_21_197

   -- array reader array_reader_198
   process(s238_0, s238_1, s238_2, s238_3, s238_4, s238_5, s238_6, s238_7, s238_8, s238_9, s238_10, s238_11, s238_12, s238_13, s238_14, s238_15, s238_16, s238_17, s238_18, s238_19, s238_20, s238_21, s238_22, s240)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s240, const00000) = '1' ) then s241 <= s238_0; else
       if (equal(s240, const00001) = '1' ) then s241 <= s238_1; else
       if (equal(s240, const00010) = '1' ) then s241 <= s238_2; else
       if (equal(s240, const00011) = '1' ) then s241 <= s238_3; else
       if (equal(s240, const00100) = '1' ) then s241 <= s238_4; else
       if (equal(s240, const00101) = '1' ) then s241 <= s238_5; else
       if (equal(s240, const00110) = '1' ) then s241 <= s238_6; else
       if (equal(s240, const00111) = '1' ) then s241 <= s238_7; else
       if (equal(s240, const01000) = '1' ) then s241 <= s238_8; else
       if (equal(s240, const01001) = '1' ) then s241 <= s238_9; else
       if (equal(s240, const01010) = '1' ) then s241 <= s238_10; else
       if (equal(s240, const01011) = '1' ) then s241 <= s238_11; else
       if (equal(s240, const01100) = '1' ) then s241 <= s238_12; else
       if (equal(s240, const01101) = '1' ) then s241 <= s238_13; else
       if (equal(s240, const01110) = '1' ) then s241 <= s238_14; else
       if (equal(s240, const01111) = '1' ) then s241 <= s238_15; else
       if (equal(s240, const10000) = '1' ) then s241 <= s238_16; else
       if (equal(s240, const10001) = '1' ) then s241 <= s238_17; else
       if (equal(s240, const10010) = '1' ) then s241 <= s238_18; else
       if (equal(s240, const10011) = '1' ) then s241 <= s238_19; else
       if (equal(s240, const10100) = '1' ) then s241 <= s238_20; else
       if (equal(s240, const10101) = '1' ) then s241 <= s238_21; else
       s241 <= s238_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_199
   process(s133, s241, s239)
   begin
   if ( s133 = '1') then s242 <= s239; else s242 <= s241;
   end if;
   end process;

   -- array writer array_writer_200
   process(s238_0, s238_1, s238_2, s238_3, s238_4, s238_5, s238_6, s238_7, s238_8, s238_9, s238_10, s238_11, s238_12, s238_13, s238_14, s238_15, s238_16, s238_17, s238_18, s238_19, s238_20, s238_21, s238_22, s240, s242)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s240, const00000) = '1' then s243_0 <= s242; else s243_0 <= s238_0; end if;
     if equal(s240, const00001) = '1' then s243_1 <= s242; else s243_1 <= s238_1; end if;
     if equal(s240, const00010) = '1' then s243_2 <= s242; else s243_2 <= s238_2; end if;
     if equal(s240, const00011) = '1' then s243_3 <= s242; else s243_3 <= s238_3; end if;
     if equal(s240, const00100) = '1' then s243_4 <= s242; else s243_4 <= s238_4; end if;
     if equal(s240, const00101) = '1' then s243_5 <= s242; else s243_5 <= s238_5; end if;
     if equal(s240, const00110) = '1' then s243_6 <= s242; else s243_6 <= s238_6; end if;
     if equal(s240, const00111) = '1' then s243_7 <= s242; else s243_7 <= s238_7; end if;
     if equal(s240, const01000) = '1' then s243_8 <= s242; else s243_8 <= s238_8; end if;
     if equal(s240, const01001) = '1' then s243_9 <= s242; else s243_9 <= s238_9; end if;
     if equal(s240, const01010) = '1' then s243_10 <= s242; else s243_10 <= s238_10; end if;
     if equal(s240, const01011) = '1' then s243_11 <= s242; else s243_11 <= s238_11; end if;
     if equal(s240, const01100) = '1' then s243_12 <= s242; else s243_12 <= s238_12; end if;
     if equal(s240, const01101) = '1' then s243_13 <= s242; else s243_13 <= s238_13; end if;
     if equal(s240, const01110) = '1' then s243_14 <= s242; else s243_14 <= s238_14; end if;
     if equal(s240, const01111) = '1' then s243_15 <= s242; else s243_15 <= s238_15; end if;
     if equal(s240, const10000) = '1' then s243_16 <= s242; else s243_16 <= s238_16; end if;
     if equal(s240, const10001) = '1' then s243_17 <= s242; else s243_17 <= s238_17; end if;
     if equal(s240, const10010) = '1' then s243_18 <= s242; else s243_18 <= s238_18; end if;
     if equal(s240, const10011) = '1' then s243_19 <= s242; else s243_19 <= s238_19; end if;
     if equal(s240, const10100) = '1' then s243_20 <= s242; else s243_20 <= s238_20; end if;
     if equal(s240, const10101) = '1' then s243_21 <= s242; else s243_21 <= s238_21; end if;
     if equal(s240, const10110) = '1' then s243_22 <= s242; else s243_22 <= s238_22; end if;
   end process;

   s245 <= "10110";  -- constint module constint_22_201

   -- array reader array_reader_202
   process(s243_0, s243_1, s243_2, s243_3, s243_4, s243_5, s243_6, s243_7, s243_8, s243_9, s243_10, s243_11, s243_12, s243_13, s243_14, s243_15, s243_16, s243_17, s243_18, s243_19, s243_20, s243_21, s243_22, s245)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
       if (equal(s245, const00000) = '1' ) then s246 <= s243_0; else
       if (equal(s245, const00001) = '1' ) then s246 <= s243_1; else
       if (equal(s245, const00010) = '1' ) then s246 <= s243_2; else
       if (equal(s245, const00011) = '1' ) then s246 <= s243_3; else
       if (equal(s245, const00100) = '1' ) then s246 <= s243_4; else
       if (equal(s245, const00101) = '1' ) then s246 <= s243_5; else
       if (equal(s245, const00110) = '1' ) then s246 <= s243_6; else
       if (equal(s245, const00111) = '1' ) then s246 <= s243_7; else
       if (equal(s245, const01000) = '1' ) then s246 <= s243_8; else
       if (equal(s245, const01001) = '1' ) then s246 <= s243_9; else
       if (equal(s245, const01010) = '1' ) then s246 <= s243_10; else
       if (equal(s245, const01011) = '1' ) then s246 <= s243_11; else
       if (equal(s245, const01100) = '1' ) then s246 <= s243_12; else
       if (equal(s245, const01101) = '1' ) then s246 <= s243_13; else
       if (equal(s245, const01110) = '1' ) then s246 <= s243_14; else
       if (equal(s245, const01111) = '1' ) then s246 <= s243_15; else
       if (equal(s245, const10000) = '1' ) then s246 <= s243_16; else
       if (equal(s245, const10001) = '1' ) then s246 <= s243_17; else
       if (equal(s245, const10010) = '1' ) then s246 <= s243_18; else
       if (equal(s245, const10011) = '1' ) then s246 <= s243_19; else
       if (equal(s245, const10100) = '1' ) then s246 <= s243_20; else
       if (equal(s245, const10101) = '1' ) then s246 <= s243_21; else
       s246 <= s243_22;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
       end if;
   end process;

   -- mux2x1 module mux2x1_203
   process(s133, s246, s244)
   begin
   if ( s133 = '1') then s247 <= s244; else s247 <= s246;
   end if;
   end process;

   -- array writer array_writer_204
   process(s243_0, s243_1, s243_2, s243_3, s243_4, s243_5, s243_6, s243_7, s243_8, s243_9, s243_10, s243_11, s243_12, s243_13, s243_14, s243_15, s243_16, s243_17, s243_18, s243_19, s243_20, s243_21, s243_22, s245, s247)
       constant const00000 : std_logic_vector(4 downto 0) := "00000";
       constant const00001 : std_logic_vector(4 downto 0) := "00001";
       constant const00010 : std_logic_vector(4 downto 0) := "00010";
       constant const00011 : std_logic_vector(4 downto 0) := "00011";
       constant const00100 : std_logic_vector(4 downto 0) := "00100";
       constant const00101 : std_logic_vector(4 downto 0) := "00101";
       constant const00110 : std_logic_vector(4 downto 0) := "00110";
       constant const00111 : std_logic_vector(4 downto 0) := "00111";
       constant const01000 : std_logic_vector(4 downto 0) := "01000";
       constant const01001 : std_logic_vector(4 downto 0) := "01001";
       constant const01010 : std_logic_vector(4 downto 0) := "01010";
       constant const01011 : std_logic_vector(4 downto 0) := "01011";
       constant const01100 : std_logic_vector(4 downto 0) := "01100";
       constant const01101 : std_logic_vector(4 downto 0) := "01101";
       constant const01110 : std_logic_vector(4 downto 0) := "01110";
       constant const01111 : std_logic_vector(4 downto 0) := "01111";
       constant const10000 : std_logic_vector(4 downto 0) := "10000";
       constant const10001 : std_logic_vector(4 downto 0) := "10001";
       constant const10010 : std_logic_vector(4 downto 0) := "10010";
       constant const10011 : std_logic_vector(4 downto 0) := "10011";
       constant const10100 : std_logic_vector(4 downto 0) := "10100";
       constant const10101 : std_logic_vector(4 downto 0) := "10101";
       constant const10110 : std_logic_vector(4 downto 0) := "10110";
   begin
     if equal(s245, const00000) = '1' then s248_0 <= s247; else s248_0 <= s243_0; end if;
     if equal(s245, const00001) = '1' then s248_1 <= s247; else s248_1 <= s243_1; end if;
     if equal(s245, const00010) = '1' then s248_2 <= s247; else s248_2 <= s243_2; end if;
     if equal(s245, const00011) = '1' then s248_3 <= s247; else s248_3 <= s243_3; end if;
     if equal(s245, const00100) = '1' then s248_4 <= s247; else s248_4 <= s243_4; end if;
     if equal(s245, const00101) = '1' then s248_5 <= s247; else s248_5 <= s243_5; end if;
     if equal(s245, const00110) = '1' then s248_6 <= s247; else s248_6 <= s243_6; end if;
     if equal(s245, const00111) = '1' then s248_7 <= s247; else s248_7 <= s243_7; end if;
     if equal(s245, const01000) = '1' then s248_8 <= s247; else s248_8 <= s243_8; end if;
     if equal(s245, const01001) = '1' then s248_9 <= s247; else s248_9 <= s243_9; end if;
     if equal(s245, const01010) = '1' then s248_10 <= s247; else s248_10 <= s243_10; end if;
     if equal(s245, const01011) = '1' then s248_11 <= s247; else s248_11 <= s243_11; end if;
     if equal(s245, const01100) = '1' then s248_12 <= s247; else s248_12 <= s243_12; end if;
     if equal(s245, const01101) = '1' then s248_13 <= s247; else s248_13 <= s243_13; end if;
     if equal(s245, const01110) = '1' then s248_14 <= s247; else s248_14 <= s243_14; end if;
     if equal(s245, const01111) = '1' then s248_15 <= s247; else s248_15 <= s243_15; end if;
     if equal(s245, const10000) = '1' then s248_16 <= s247; else s248_16 <= s243_16; end if;
     if equal(s245, const10001) = '1' then s248_17 <= s247; else s248_17 <= s243_17; end if;
     if equal(s245, const10010) = '1' then s248_18 <= s247; else s248_18 <= s243_18; end if;
     if equal(s245, const10011) = '1' then s248_19 <= s247; else s248_19 <= s243_19; end if;
     if equal(s245, const10100) = '1' then s248_20 <= s247; else s248_20 <= s243_20; end if;
     if equal(s245, const10101) = '1' then s248_21 <= s247; else s248_21 <= s243_21; end if;
     if equal(s245, const10110) = '1' then s248_22 <= s247; else s248_22 <= s243_22; end if;
   end process;

   s249 <= '0';  -- constint module constint_0_205

   -- mux2x1 module mux2x1_206
   process(s133, s128, s249)
   begin
   if ( s133 = '1') then s250 <= s249; else s250 <= s128;
   end if;
   end process;

   s251 <= s131 or s133;  -- or2 or2_207

   s252 <= s40 or s251;  -- or2 or2_208

   -- register state_reg_209
   process (s3, s4, s5)
   begin
   if s5 = '1' then
     s253 <= '0';
   elsif s3'event and s3='1' then  
     if s4 = '1' then
        s253 <= '0';
     else
        s253 <= s252;
     end if;
   end if;
   end process;

   s7 <= s6 or s253;  -- or2 or2_210

   s9 <= s7 and s8;  -- and2 and2_211

   s256 <= not s8;  -- not module inv_212

   s257 <= s7 and s256;  -- and2 and2_213

   s302 <= '0';  -- constint module constint_0_224

   s303 <= '1';  -- constint module constint_minus1_225

   s306 <= "11111";  -- constint module constint_31_226

   -- bitselect bitselect_227
   s305 <= s57(to_integer(to_unsigned(s306)));

   -- mux2x1 module mux2x1_228
   process(s305, s302, s303)
   begin
   if ( s305 = '1') then s304 <= s303; else s304 <= s302;
   end if;
   end process;

   s59 <= s304 & s57;  -- concat module concat_module_229

   s309 <= '0';  -- constint module constint_0_231

   s310 <= '1';  -- constint module constint_minus1_232

   s313 <= "11111";  -- constint module constint_31_233

   -- bitselect bitselect_234
   s312 <= s63(to_integer(to_unsigned(s313)));

   -- mux2x1 module mux2x1_235
   process(s312, s309, s310)
   begin
   if ( s312 = '1') then s311 <= s310; else s311 <= s309;
   end if;
   end process;

   s68 <= s311 & s63;  -- concat module concat_module_236

   s316 <= "00000000000000000000000000000";  -- constint module constint_0_238

   s317 <= "11111111111111111111111111111";  -- constint module constint_minus1_239

   s320 <= "100011";  -- constint module constint_35_240

   -- bitselect bitselect_241
   s319 <= s91(to_integer(to_unsigned(s320)));

   -- mux2x1 module mux2x1_242
   process(s319, s316, s317)
   begin
   if ( s319 = '1') then s318 <= s317; else s318 <= s316;
   end if;
   end process;

   s103 <= s318 & s91;  -- concat module concat_module_243

   s323 <= "0000000000000000000000000000000000000000000000";  -- constint module constint_0_245

   s324 <= "1111111111111111111111111111111111111111111111";  -- constint module constint_minus1_246

   s327 <= "10001";  -- constint module constint_17_247

   -- bitselect bitselect_248
   s326 <= s106(to_integer(to_unsigned(s327)));

   -- mux2x1 module mux2x1_249
   process(s326, s323, s324)
   begin
   if ( s326 = '1') then s325 <= s324; else s325 <= s323;
   end if;
   end process;

   s107 <= s325 & s106;  -- concat module concat_module_250

   s330 <= "00000000000000000000000000000000";  -- constint module constint_0_252

   s331 <= "11111111111111111111111111111111";  -- constint module constint_minus1_253

   s334 <= "11111";  -- constint module constint_31_254

   -- bitselect bitselect_255
   s333 <= s110(to_integer(to_unsigned(s334)));

   -- mux2x1 module mux2x1_256
   process(s333, s330, s331)
   begin
   if ( s333 = '1') then s332 <= s331; else s332 <= s330;
   end if;
   end process;

   s111 <= s332 & s110;  -- concat module concat_module_257

   s337 <= '0';  -- constint module constint_0_259

   s338 <= '1';  -- constint module constint_minus1_260

   s341 <= "111111";  -- constint module constint_63_261

   -- bitselect bitselect_262
   s340 <= s112(to_integer(to_unsigned(s341)));

   -- mux2x1 module mux2x1_263
   process(s340, s337, s338)
   begin
   if ( s340 = '1') then s339 <= s338; else s339 <= s337;
   end if;
   end process;

   s113 <= s339 & s112;  -- concat module concat_module_264
end SynFir_DoCalculate_syn;

